--------------------------------------------------------------------------------
-- Company:        vienna university of technology
-- Engineer:       mario faschang
-- Create Date:    11:12:56 19/01/2010
-- Module Name:    tb_ClkGen
-- Project Name:   i2c master controller
-- Description:  * testbench for the variable Clock-Generator
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
USE ieee.numeric_std.ALL;

ENTITY tb_ClkDiv IS
END tb_ClkDiv;

