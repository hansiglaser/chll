--------------------------------------------------------------------------------
-- Company:        vienna university of technology
-- Engineer:       mario faschang
-- Create Date:    11:12:56 19/01/2010
-- Module Name:    tb_I2CTransferController
-- Project Name:   i2c master controller
-- Description:  * testbench for i2cTransferController
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY tb_I2CTransferController IS
END tb_I2CTransferController;

