package Config is

  constant CfgClkGating : boolean := false;

end Config;

package body Config is

end Config;
