  constant TRFSM1Length : integer := 1778;
  constant TRFSM1Cfg    : std_logic_vector(TRFSM1Length-1 downto 0) := "00000100011100001001100100000010000000000000011100000000010100101000000100101000000011000001100000100100001000011100010000001001100010000100000010100000100101000000100100001000001000010000011111100000000000000000000011111100000000000000000000011111100000000000000000000000000000000001000100000000000011100000000000000000001001000011000000100100000000001000000000010100001000000001010000100001000000000011000100000000100100000100001100000000101000001100000000100000000001100000000100100100100001000100000000101000000000100100000100001000100000000101000000000101000101000000000100000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000000111111000000000000000000000000000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000111111000000000000000000000000000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000";
