  constant SensorFSMLength : integer := 850;
  constant SensorFSMCfg    : std_logic_vector(SensorFSMLength-1 downto 0) := "0010000011000001010011111000000000000000111110000000000000001111100000000000000011111000000000000000000000000000001010000000000100000000000000000011000011000000100000001000000000101000000000010000000010000000001100000100000100000001000000001001000001000001010000010000000011000010001000000100000001100000000010101000000000001000000110000001001100000010000000100100011000000100100100001100000010001111100000000000000000000000000000000100000100110001000000001100000100001111100000000000000000000000000000000011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000000010000011011000000000000000100001100000100000001000001101100000000000100000001000000001010111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
