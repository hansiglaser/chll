--------------------------------------------------------------------------------
-- Company:        vienna university of technology
-- Engineer:       mario faschang
-- Create Date:    11:22:56 11/26/2009
-- Module Name:    tb_I2CCore
-- Project Name:   i2c master controller
-- Description:  * testbench for i2ccore
--               * generates different scenarios of the i2c-bus-communication
--                 to verify the behavior of the i2c-core.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY tb_I2CCore IS
END tb_I2CCore;

