

architecture structure of RxModule is

-- signal declaration

  -- signals for Rx module
  signal SamplingBaudClk            : std_logic;
  signal RxParityError              : std_logic;
  signal RxStopBitError             : std_logic;
  signal RxBufferFullError          : std_logic;
  signal RxFifoFull                 : std_logic;
  signal RxBGEnable                 : std_logic;
  signal RxStateMachineParallelData : std_logic_vector((MaxDataWidth-1) downto 0);
  signal RxSaveData                 : std_logic;
  signal RxBaudClk                  : std_logic;

-- component declaration

  component BaudGenerator
    generic ( MaxSpeedDividerWidth : integer);
    Port    ( Clk_i                : in  STD_LOGIC;
              Reset_i_n            : in  STD_LOGIC;
              BGEnable_i           : in  STD_LOGIC;
              SpeedDivider_i       : in  STD_LOGIC_VECTOR((MaxSpeedDividerWidth-1) downto 0);
              BaudClk_o            : out STD_LOGIC;
              BaudSamplingClk_o    : out STD_LOGIC);
  end component;

  component RxDataStateMachine
    generic ( MaxDataWidth     : integer range 2 to 64;
              Oversampling     : integer range 2 to 3);
    Port ( Reset_i_n           : in  STD_LOGIC;
           Clk_i               : in  STD_LOGIC;
           SamplingBaudClk_i   : in  STD_LOGIC;
           BaudClk_i           : in  STD_LOGIC;
           FifoFull_i          : in  STD_LOGIC;
           BitSelect_i         : in  BitSelectionType;
           ParityOn_i          : in  STD_LOGIC;
           ParityEvenOdd_i     : in  ParityType;
           RxD_i               : in  STD_LOGIC;
           BGEnable_o          : out STD_LOGIC;
           ParallelData_o      : out STD_LOGIC_VECTOR((MaxDataWidth-1) downto 0);
           WriteParallelData_o : out STD_LOGIC;
           ParityError_o       : out STD_LOGIC;
           StopBitError_o      : out STD_LOGIC;
           RxBufferFullError_o : out STD_LOGIC);
  end component;

  component ErrorIndicator
    Port ( -- Errors generated by the TX/RX module
           ParityError_i                : in   STD_LOGIC;
           StopBitError_i               : in   STD_LOGIC;
           RxBufferFullError_i          : in   STD_LOGIC;
           -- general inputs
           Clk_i                        : in   STD_LOGIC;
           ErrorReset_i                 : in   STD_LOGIC;
           Reset_i_n                    : in   STD_LOGIC;
           -- Indication
           StopBitErrorIndicator_o      : out  STD_LOGIC;
           ParityErrorIndicator_o       : out  STD_LOGIC;
           RxBufferFullErrorIndicator_o : out  STD_LOGIC
          );
  end component;

  component FIFOSyncTop
    Generic ( DataWidth   : integer range 2 to 64;
              AdressWidth : integer range 2 to 10);
    Port    ( Reset_n     : in  STD_LOGIC;
              Clk         : in  STD_LOGIC;
              DataA_i     : in  STD_LOGIC_VECTOR (DataWidth - 1 downto 0);
              WriteA_i    : in  STD_LOGIC;
              DataB_o     : out STD_LOGIC_VECTOR (DataWidth - 1 downto 0);
              ReadNextB_i : in  STD_LOGIC;
              FIFOFull_o  : out STD_LOGIC;
              FIFOEmpty_o : out STD_LOGIC);
  end component;

begin

  -- Rx BaudGenerator
  RXBAUD: BaudGenerator
    generic map ( MaxSpeedDividerWidth => MaxSpeedDividerWidth)
    port map    ( Clk_i                => Clk_i,
                  Reset_i_n            => Reset_i_n,
                  BGEnable_i           => RxBGEnable,
                  SpeedDivider_i       => SpeedDivider_i,
                  BaudClk_o            => RxBaudClk,
                  BaudSamplingClk_o    => SamplingBaudClk);

  -- RxDataStateMachine
  RXSM: RxDataStateMachine
    generic map ( MaxDataWidth        => MaxDataWidth,
                  Oversampling        => Oversampling)
    port map    ( Reset_i_n           => Reset_i_n,
                  Clk_i               => Clk_i,
                  SamplingBaudClk_i   => SamplingBaudClk,
                  BaudClk_i           => RxBaudClk,
                  FifoFull_i          => RxFifoFull,
                  BitSelect_i         => BitsSelect_i,
                  ParityOn_i          => ParityOn_i,
                  ParityEvenOdd_i     => ParityEvenOdd_i,
                  RxD_i               => RxD_i,
                  BGEnable_o          => RxBGEnable,
                  ParallelData_o      => RxStateMachineParallelData,
                  WriteParallelData_o => RxSaveData,
                  ParityError_o       => RxParityError,
                  StopBitError_o      => RxStopBitError,
                  RxBufferFullError_o => RxBufferFullError);

  -- Rx ErrorIndicator
  RXERRORIND: ErrorIndicator
    port map    ( -- Errors generated by the TX/RX module
                  ParityError_i                 => RxParityError,
                  StopBitError_i                => RxStopBitError,
                  RxBufferFullError_i           => RxBufferFullError,
                  -- general inputs
                  Clk_i                         => Clk_i,
                  ErrorReset_i                  => ErrorReset_i,
                  Reset_i_n                     => Reset_i_n,
                  -- Indication
                  StopBitErrorIndicator_o       => RxStopBitErrorIndicator_o,
                  ParityErrorIndicator_o        => RxParityErrorIndicator_o,
                  RxBufferFullErrorIndicator_o  => RxBufferFullErrorIndicator_o);

  -- Rx Fifo
  RXFIFO: FIFOSyncTop
    generic map ( DataWidth   => MaxDataWidth,
                  AdressWidth => RxFifoAdressWidth)
    port map    ( Reset_n     => Reset_i_n,
                  Clk         => Clk_i,
                  DataA_i     => RxStateMachineParallelData,
                  WriteA_i    => RxSaveData,
                  DataB_o     => RxData_o,
                  ReadNextB_i => RxRd_i,
                  FIFOFull_o  => RxFifoFull,
                  FIFOEmpty_o => RxEmpty_o);

  RxFull_o  <= RxFifoFull;

end structure;

