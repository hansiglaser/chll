  constant SensorFSMLength : integer := 850;
  constant SensorFSMCfg    : std_logic_vector(SensorFSMLength-1 downto 0) := "0001100010000000000011111000000000000000111110000000000000001111100000000000000011111000000000000000000000000000001010000000000000100000000000000011000010000000001000001000000001001000010000000100000100000000001010000000000000011111100000000000000000000000000000001000000011000100001000000001000000100000001101000000110000000100000100000001001100000001000000000100010000000100100100001000000000011111100000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
