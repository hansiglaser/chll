  constant FSMLength : integer := 1295;
  constant FSMCfg    : std_logic_vector(FSMLength-1 downto 0) := "00010001010000000010100100010000011000000001000001111110000000000000000000011111000000000000000000001111100000000000000000000000000000001001000000000000010000000000000000010100001100000000010000000001000000010100001000000001011010000110000001001000000000000010000000010100000100100000100000000101101000101000001000100101000000001010010111110000000000000000000000000000001111100000000000000000000000000000011111000000000000000000000000000000111110000000000000000000000000000000000100100001100000011000000001011010000110000101010000001000000000101000000011000010100010000110000000001000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000000010011000100000010000110000000010110100000100110001000010000010000000000101111011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
