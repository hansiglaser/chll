  constant bitdataLength : integer := 1282;
  constant bitdataCfg    : std_logic_vector(bitdataLength-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000101011010100000000000000100100000000100000000000000000000000000000000001000000000000000000000000000000000010001000001000000000000110010010000110000000000010001011000000000000000000000000000100100000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101010110110100000110010000000000000000000000000100110101011100000000000011110100101010001000010001010001001100000000000000000000000000000000000000000100011001000110001100011000110011101011000000100001111011010100011000110001100010000011000010001101000000010001111011010100010000111000001001010001010000000000000000000001000000000011000001110101000000000000010000010100010110100000000000000000000000100000001000100000000011010100010100000010000011100011001101011000000000000001100101000000000001000100000000000000000000000000001000000000000000000000000000000001001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000";
