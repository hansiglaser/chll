  constant SensorFSMLength : integer := 850;
  constant SensorFSMCfg    : std_logic_vector(SensorFSMLength-1 downto 0) := "0001100010000001100011111000000000000000111110000000000000001111100000000000000011111000000000000000000000000000001010000000000010000000000000000011000010000000010000001000000001001000010000001000000100000000001010000000000001001111100000000000000000000000000000001000001001010000001000000010000001000000001011000000010000000101000100000000101001000010000000010011111000000000000000000000000000001111100000000000000000000000000000000010000011010000000100001000000010000000100000110100000100000011000000011011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
