  constant FSMLength : integer := 1295;
  constant FSMCfg    : std_logic_vector(FSMLength-1 downto 0) := "00010001010000000000001000010000011000000000100000111110000000000000000000011111000000000000000000001111100000000000000000000000000000010001000000000000000100000000000000100100001100000000001000000001000000010100001000000000000001000110000010001000000000000000010000010100001000100000100000000000001000101000010000100101000000000000010111110000000000000000000000000000001111100000000000000000000000000000011111000000000000000000000000000000111110000000000000000000000000000000000100000011001000011000000000000001000010000001110000010000000000000000100011000101001000000100000000000010000001100010100001000011000000000001000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
