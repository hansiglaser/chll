  constant TRFSM0Length : integer := 820;
  constant TRFSM0Cfg    : std_logic_vector(TRFSM0Length-1 downto 0) := "0000100100000000101000010001010000000000000110001000000100001111100000000000000011111000000000000000111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000000000000001010000000001000000000000000110000110000010000001000000010100000000010000100100000001100001100000100010010100001001000010000001100001010000101000101000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000001111100000000000000000000000001111100000000000000000000000001111100000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000000000000111110000000000000000000000000000000000000";
