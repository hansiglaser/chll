----------------------------------------------------------------------------------
-- Company:     TU Vienna
-- Engineer:    Georg Blemenschitz
--
-- Create Date: 20:52:31 01/31/2010
-- Design Name: SPI
-- Module Name: tb_SPIShifter
-- Description: VHDL Test Bench for module: SPIShifter
--
-- Revision:
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_SPIShifter is
end tb_SPIShifter;

