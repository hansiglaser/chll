  constant I2CFSMLength : integer := 1295;
  constant I2CFSMCfg    : std_logic_vector(I2CFSMLength-1 downto 0) := "00011000000001000000000000010001010000000100000000001100110000000000001000000111001000000010000000000100000101000000000000010000000000100001000000000100000000000000000001000100011100001000000000000001000000011000001000000000000100000010000000101010000000000000001000001000000010100000000000000100000000101000000011000101000000000000001001010000000101010110000000000000010100100000100100011000000000010000001001000001000101001000000000100000010100000000011000100000000100000000001000000011001000010000000001000000000100000001100010100100000000100000001011000000001111000110010000000000000110000000000111100001000000000001000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
