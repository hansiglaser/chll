  constant TRFSM0Length : integer := 820;
  constant TRFSM0Cfg    : std_logic_vector(TRFSM0Length-1 downto 0) := "0010000011000001010011111000000000000000111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000000000000001010000000000100000000000000110000110000001000000010000010100000000001000000001000001100000100000100000001000010010000010000010100000110000010100000000000100011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000000001000011000010001000000100000001100100110000001000000010010001100100100100001100000010001111100000000000000000000000000001010011000100000000110000010000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000000101101100000000000000010000110000010000000101101100000000000100000001000000001010";
