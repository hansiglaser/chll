  constant TRFSM1Length : integer := 1778;
  constant TRFSM1Cfg    : std_logic_vector(TRFSM1Length-1 downto 0) := "00000100010100000000000100100001000011000000000000000000001100000000000000001001000010000001000000000010000000010100001100000000001001011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000000000000000000010100000000000000001000000000000000000011000010000000000010000000011000000000100100000100000000000110000011000000000101000011000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000000111111000000000000000000000000000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000111111000000000000000000000000000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000";
