----------------------------------------------------------------------------------
-- Company:     TU Vienna
-- Engineer:    Georg Blemenschitz
-- 
-- Create Date: 17:41:00 01/18/2010 
-- Design Name: SPI
-- Module Name: tb_SPI 
-- Description: VHDL Test Bench for module: SPI
--
-- Revision: 
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
 
entity tb_SPI is
end tb_SPI;

