  constant bitdataLength : integer := 1282;
  constant bitdataCfg    : std_logic_vector(bitdataLength-1 downto 0) := "0000000000000000001000001001000010010001000000110000001000000000100000000000000000000011000011000000000000000000000000000000000000000001000000000000000000000000000000000010001000100000000000000000000000000000000000000010000000011000000000000000000000001001000000010000001000000000000000000000000000000000000000000001001000001000100011010000100100001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101000000000000000001110000000000001000000000000000101100000000000000000101001101110110000010000101000000011010110101101011010110101101010000001100000000000000000000000000100100010000000111100100000000000000000000000000000000001101101011100100110000000000000000000000000000000000000000000000000000000000000000000000000110100000110000100011010100000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000111000100010101100000000000000000000000101100000011110000101110000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110001000000000011100000000000000000001010010000001001000000000000000010000100000001010000000000000000000000000000000000000000000000000000000000000000000000000000";
