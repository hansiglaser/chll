  constant bitdataLength : integer := 1282;
  constant bitdataCfg    : std_logic_vector(bitdataLength-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000101011010100000000000000100000100000000000000001100000011000000000000011000000000000000000000000000000000010001000100000000000000000000000000000000000000000000011000000000000000000000000000100100000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110110100000000000000000000000000000000000000110101011101001010100010000000000000000000000000000110001100000000000000000000000000000000000000000100011001000110001100011000110001100011000110001101101010000100010000000000010010100000000110100100000000000000000000000000000011011000010001111001110000000000000000000000000000000001000000000000000000000000000000011000100110100000000000000000000001000000010000000000000000000000010100000000000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001011000000000011100000000000000000000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
