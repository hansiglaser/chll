  constant TRFSM2Length : integer := 1020;
  constant TRFSM2Cfg    : std_logic_vector(TRFSM2Length-1 downto 0) := "001000001100000101001111100000000000000011111000000000000000111110000000000000001111100000000000000000000000000000101000000000010000000000000000001100001100000010000000100000000010100000000001000000001000000000110000010000010000000100000000100100000100000101000001000000001100001000100000010000000110000000001010100000000000100000011000000100110000001000000010010001100000010010010000110000001000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000000100000100110001000000001100000100001111100000000000000000000000000000000011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000000010000011011000000000000000100001100000100000001000001101100000000000100000001000000001010111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
