  constant TRFSM0Length : integer := 820;
  constant TRFSM0Cfg    : std_logic_vector(TRFSM0Length-1 downto 0) := "0001000101000101001000100000110001000001111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000000000000010010000000010000000000000001010000110000100000000010000010100001000101101000011000010010000000010000000010100010010000010001011010001010001000100101000101001011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000000000110000110000001100010110100001100101010000001000010100000001100101000100001100001000001111100000000000000000000000000000111000100000010000110001011010000011100010000100000100000101111011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000000000000111110000000000000000000000000000000000000";
