  constant SensorFSMLength : integer := 850;
  constant SensorFSMCfg    : std_logic_vector(SensorFSMLength-1 downto 0) := "0010000011000000000111111000000000000000111110000000000000001111100000000000000011111000000000000000000000000000001010000000000010000000000000000011000011000000100000001000000000101000000000000000000010000000001100000100000000000001000000001001000001000000001000010000000011000010001000000000100001100000000010101000000000000100000110000010001100000010000000010000011000001000100100001100000001001111100000000000000000000000000000000100000001110000000100001100000000100001000000011100010000000100000000001011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
