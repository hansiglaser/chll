  constant TRFSM0Length : integer := 820;
  constant TRFSM0Cfg    : std_logic_vector(TRFSM0Length-1 downto 0) := "0001100010000001100011111000000000000000111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000000000000001010000000000010000000000000110000100000000100000010000100100001000000100000010000001010000000000001001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000000000101001010000001000000010000001000010110000000100000001010001000010100100001000000001001111100000000000000000000000000000101101000000010000100000001000000010110100000100000011000000011011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000000000000111110000000000000000000000000000000000000";
