----------------------------------------------------------------------------------
-- Company:     TU Vienna
-- Engineer:    Georg Blemenschitz
--
-- Create Date: 09:33:07 01/29/2010
-- Design Name: SPI
-- Module Name: tb_SPIControl
-- Description: VHDL Test Bench for module: SPIControl
--
-- Revision:
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_SPIControl is
end tb_SPIControl;

