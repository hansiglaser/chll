  constant SPIFSMLength : integer := 1295;
  constant SPIFSMCfg    : std_logic_vector(SPIFSMLength-1 downto 0) := "00001001110000010000000000010000000000000000000000001010101000000000100000000110000110000000000010000011100100000000100000000000000000010001000000000000000100000000000000100100011000000000001000000010000000010100010000000000000001000100000000110010000000000000000010001100000010100001100000000000010000011000000100101001000000000000100010000000000011001010000000100000000100100000000110001000000000000001001010000000100100001000000000100000010100000001010010100000000001000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
