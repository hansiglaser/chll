  constant bitdataLength : integer := 1282;
  constant bitdataCfg    : std_logic_vector(bitdataLength-1 downto 0) := "0000000000000000001000000101000011111111000000000000000000001000100000000000000000000011000011000000000000000000000000000000000000000001000000000000000000000000000000000010001000100000000000000000000000000000000000000010001011000000000000000000000000000100100000000000001000011000000000000000000000000100000000000001001000000000000000000000000100001000001000000000000000000000000000000000000000000000000000000001110110100000000000000000000000000000000000000110101011100000000000011110000000000001000000000000000101100000000000000000000000000000000000000000100011001000110001100011000110001100011000110100001101000000100010000000000000001001000000101100100000000000000000000000000000000000000101101100110001000000000000000000000000001010001000000000000000000000000000000000000000110100000000000000000000010000000010000000000000000000000000100000000000000000000000000011010011100000000000001000000000000000000000000000000000000000000000000000001000100110001110000000011001110000000000000000000000000000011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001011000100000011100000000000000001110000010000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
