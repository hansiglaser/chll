  constant SensorFSMLength : integer := 1180;
  constant SensorFSMCfg    : std_logic_vector(SensorFSMLength-1 downto 0) := "0011000101100000000011111000000000000000111110000000000000001111100000000000000011111000000000000000000000000000001010000000000001000000000000000011000101000000010000001000000010001000010100000000000010000000100100011001000000000001000000001000100010000001000000010000000010010001110000010000000110000000100010001100000000010001100000001001001000000000000100100000000010001001000001000000001000000000100100100100010000000010100000000010101000000000000010001010000001001100000011000000001000101000000100100100010100000000100011100000000101100001000000100000001110000000010001100111000010000001000000000001011000001000000010000100000000000100011010000000001000010010000000010110000001001000000001001000000001000110100100100000001111100000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
