  constant TRFSM1Length : integer := 1778;
  constant TRFSM1Cfg    : std_logic_vector(TRFSM1Length-1 downto 0) := "11111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000000000000000000010100000000000001001000000000000000000011000010100000001000100000000100000001000100000100000001001000000000100000001001000011000000001011000000001000000001000100001000000001001000000001000000001001000011100000000111000000001100000001000100001100000001001000000001100000001001000100000000000111001000010000000001000100010000000001001000000010000000001001000100100000000111000000010100000000010100000000000001000100000011000001000001000010100000001001000000011100000000101000010000000000101010000011100000000100100011100000000101000000100000000000101000001000000000101010000100000000000100100100000000000101000000100100000000101000000100000000101010000100100000000100100100100000000101000011111100000000000000000000000000000000011111100000000000000000000000000000000000010100000010011000000011000000010001100000101000000100100100001010000000100010000001100000110000000100010100000001001000000011000001100000010000101000000010010001111111000000000000000000000000000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000";
