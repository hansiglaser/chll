  constant I2CFSMLength : integer := 1295;
  constant I2CFSMCfg    : std_logic_vector(I2CFSMLength-1 downto 0) := "00011000000010000000010000010001010011000000000010001100110001100000000000000111001000110000000001000100000101001000001100000000000000100001000000010000100000000000000001000100011101100001000000000001000000011000001001000000000001000010000000101010000110000000000010001000000010100000000100010000000000101000000011000101001000000100000001010000000101010110010110001000000100100000100100011001100001000000001001000001000101001000100010000000010100000000011000100010000010000000001000000011001000010001000000000000000100000001100010100100010000000000001011000000001111000110010100000100000110000000000111100001001000001000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
