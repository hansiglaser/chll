  constant TRFSM2Length : integer := 1020;
  constant TRFSM2Cfg    : std_logic_vector(TRFSM2Length-1 downto 0) := "000010010000000010100001000101000000000000011000100000010000111110000000000000001111100000000000000000000000000000101000000000100000000000000000001100001100000100000010000000000010100000000010000100100000000000110000110000010001001010000000010010000100000011000010100000000101100001010000000000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000011111000000000000000000000000000001111100000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
