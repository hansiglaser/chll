configuration MyReconfigLogicTestParamIntf_cfg of MyReconfigLogic is
  for TestParamIntf
  end for;
end MyReconfigLogicTestParamIntf_cfg;
