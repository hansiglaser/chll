  constant bitdataLength : integer := 1282;
  constant bitdataCfg    : std_logic_vector(bitdataLength-1 downto 0) := "0000000000000000001000001001000010010001000000110000001000000000100000000000000000000011000011000000000000000000000000011000000000000011000000000000000000000000000000000010001000100000010110000000000000000000000000000000000011000000000000000000000000001001000000010000001000000000000000000000000000000000000000000001001000001000100011010000100100001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101011100000000000010000000000000000000000000000000101101010000000001100000000000000000000011000101000000011010110101101011010110101101010000000000000000000000000000010001100100010000000111100100000000000000000000000000000000000000000001100100110000000000000000000000000000000000000000000000000000000000000000000000000110100000000000000011010100000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000001000111000100010101100000000001101011000000101100000011110000101110000001011000000000000000000000000000000000000000000000000000000000000000000000011010000000000000000000000000000010010110000000000000011100000000000000000000000000000001001000000101100100010000100000001010000000000000000000000000000000000000010000000000000000000000000000000000000";
