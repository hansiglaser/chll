  constant SensorFSMLength : integer := 1180;
  constant SensorFSMCfg    : std_logic_vector(SensorFSMLength-1 downto 0) := "1111100000000000000011111000000000000000111110000000000000001111100000000000000011111000000000000000000000000000001010000000100100000000000000000011000101001000100000001000000010001000010010010000000010000000100100011000101100000001000000001000100010001001000000010000000010010001110001110000000110000000100010001100100100000001100000001001001000000111001000100000000010001001000010010000001000000000100100100100011100000010100000000010101000000010001000001010000001001100000011001000110000101000000100100100010100100010000011000001100000001001010010010000001100000100000110000101001001000000110000011000000100010100100100010011100000000101100001000001010100001110000000010001100111000101000001000000000001011000001000010101000100000000000100011010000001010000010010000000010110011000000100010101000100100000000100011001101001000101000011111000000000000000000000000000000000111110000000000000000000000000000000001111100000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000000000000000000000000000000000000000001111100000000000000000000000000000000000000000";
