package Config is

  constant CfgClkGating : boolean := true;

end Config;

package body Config is

end Config;
