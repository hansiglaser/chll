configuration MyReconfigLogicTestCfgIntf_cfg of MyReconfigLogic is
  for TestCfgIntf
  end for;
end MyReconfigLogicTestCfgIntf_cfg;
