module MyInterSynthModule(bitdata, AdcConvComplete_i, AdcDoConvert_o, AdcValue_i, I2C_Busy_i, I2C_DataIn_o, I2C_DataOut_i, I2C_Error_i, I2C_FIFOEmpty_i, I2C_FIFOFull_i, I2C_FIFOReadNext_o, I2C_FIFOWrite_o, I2C_ReadCount_o, I2C_ReceiveSend_n_o, I2C_StartProcess_o, Inputs_i_0, Inputs_i_1, Inputs_i_2, Inputs_i_3, Inputs_i_4, Inputs_i_5, Inputs_i_6, Inputs_i_7, Outputs_o_0, Outputs_o_1, Outputs_o_2, Outputs_o_3, Outputs_o_4, Outputs_o_5, Outputs_o_6, Outputs_o_7, ReconfModuleIRQs_o_0, ReconfModuleIRQs_o_1, ReconfModuleIRQs_o_2, ReconfModuleIRQs_o_3, ReconfModuleIRQs_o_4, SPI_CPHA_o, SPI_CPOL_o, SPI_DataIn_o, SPI_DataOut_i, SPI_FIFOEmpty_i, SPI_FIFOFull_i, SPI_LSBFE_o, SPI_ReadNext_o, SPI_Transmission_i, SPI_Write_o, ReconfModuleIn_i_0, ReconfModuleIn_i_1, ReconfModuleIn_i_2, ReconfModuleIn_i_3, ReconfModuleIn_i_4, ReconfModuleIn_i_5, ReconfModuleIn_i_6, ReconfModuleIn_i_7, ReconfModuleOut_o_0, ReconfModuleOut_o_1, ReconfModuleOut_o_2, ReconfModuleOut_o_3, ReconfModuleOut_o_4, ReconfModuleOut_o_5, ReconfModuleOut_o_6, ReconfModuleOut_o_7, ParamIn_Word_i, ParamOut_Word_o, Clk_i, Reset_n_i, CfgMode_i, CfgClk_TRFSM0_i, CfgClk_TRFSM1_i, CfgShift_TRFSM0_i, CfgShift_TRFSM1_i, CfgDataIn_i, CfgDataOut_TRFSM0_o, CfgDataOut_TRFSM1_o);

input [1281:0] bitdata;

// user inputs and outputs
input AdcConvComplete_i;
output AdcDoConvert_o;
input [15:0] AdcValue_i;
input I2C_Busy_i;
output [7:0] I2C_DataIn_o;
input [7:0] I2C_DataOut_i;
input I2C_Error_i;
input I2C_FIFOEmpty_i;
input I2C_FIFOFull_i;
output I2C_FIFOReadNext_o;
output I2C_FIFOWrite_o;
output [7:0] I2C_ReadCount_o;
output I2C_ReceiveSend_n_o;
output I2C_StartProcess_o;
input Inputs_i_0;
input Inputs_i_1;
input Inputs_i_2;
input Inputs_i_3;
input Inputs_i_4;
input Inputs_i_5;
input Inputs_i_6;
input Inputs_i_7;
output Outputs_o_0;
output Outputs_o_1;
output Outputs_o_2;
output Outputs_o_3;
output Outputs_o_4;
output Outputs_o_5;
output Outputs_o_6;
output Outputs_o_7;
output ReconfModuleIRQs_o_0;
output ReconfModuleIRQs_o_1;
output ReconfModuleIRQs_o_2;
output ReconfModuleIRQs_o_3;
output ReconfModuleIRQs_o_4;
output SPI_CPHA_o;
output SPI_CPOL_o;
output [7:0] SPI_DataIn_o;
input [7:0] SPI_DataOut_i;
input SPI_FIFOEmpty_i;
input SPI_FIFOFull_i;
output SPI_LSBFE_o;
output SPI_ReadNext_o;
input SPI_Transmission_i;
output SPI_Write_o;
input ReconfModuleIn_i_0;
input ReconfModuleIn_i_1;
input ReconfModuleIn_i_2;
input ReconfModuleIn_i_3;
input ReconfModuleIn_i_4;
input ReconfModuleIn_i_5;
input ReconfModuleIn_i_6;
input ReconfModuleIn_i_7;
output ReconfModuleOut_o_0;
output ReconfModuleOut_o_1;
output ReconfModuleOut_o_2;
output ReconfModuleOut_o_3;
output ReconfModuleOut_o_4;
output ReconfModuleOut_o_5;
output ReconfModuleOut_o_6;
output ReconfModuleOut_o_7;
input [79:0] ParamIn_Word_i;
output [31:0] ParamOut_Word_o;
input Clk_i;
input Reset_n_i;
input CfgMode_i;
input CfgClk_TRFSM0_i;
input CfgClk_TRFSM1_i;
input CfgShift_TRFSM0_i;
input CfgShift_TRFSM1_i;
input CfgDataIn_i;
output CfgDataOut_TRFSM0_o;
output CfgDataOut_TRFSM1_o;

// CellInAdcConvComplete_i[0]
wire cell_0_0; // PORT

// CellOutAdcDoConvert_o[0]
wire cell_1_0; // PORT

// CellInAdcValue_i[0]
wire [15:0] cell_2_0; // PORT

// CellInI2C_Busy_i[0]
wire cell_3_0; // PORT

// CellOutI2C_DataIn_o[0]
wire [7:0] cell_4_0; // PORT

// CellInI2C_DataOut_i[0]
wire [7:0] cell_5_0; // PORT

// CellInI2C_Error_i[0]
wire cell_6_0; // PORT

// CellInI2C_FIFOEmpty_i[0]
wire cell_7_0; // PORT

// CellInI2C_FIFOFull_i[0]
wire cell_8_0; // PORT

// CellOutI2C_FIFOReadNext_o[0]
wire cell_9_0; // PORT

// CellOutI2C_FIFOWrite_o[0]
wire cell_10_0; // PORT

// CellOutI2C_ReadCount_o[0]
wire [7:0] cell_11_0; // PORT

// CellOutI2C_ReceiveSend_n_o[0]
wire cell_12_0; // PORT

// CellOutI2C_StartProcess_o[0]
wire cell_13_0; // PORT

// CellInInputs_i_0[0]
wire cell_14_0; // PORT

// CellInInputs_i_1[0]
wire cell_15_0; // PORT

// CellInInputs_i_2[0]
wire cell_16_0; // PORT

// CellInInputs_i_3[0]
wire cell_17_0; // PORT

// CellInInputs_i_4[0]
wire cell_18_0; // PORT

// CellInInputs_i_5[0]
wire cell_19_0; // PORT

// CellInInputs_i_6[0]
wire cell_20_0; // PORT

// CellInInputs_i_7[0]
wire cell_21_0; // PORT

// CellOutOutputs_o_0[0]
wire cell_22_0; // PORT

// CellOutOutputs_o_1[0]
wire cell_23_0; // PORT

// CellOutOutputs_o_2[0]
wire cell_24_0; // PORT

// CellOutOutputs_o_3[0]
wire cell_25_0; // PORT

// CellOutOutputs_o_4[0]
wire cell_26_0; // PORT

// CellOutOutputs_o_5[0]
wire cell_27_0; // PORT

// CellOutOutputs_o_6[0]
wire cell_28_0; // PORT

// CellOutOutputs_o_7[0]
wire cell_29_0; // PORT

// CellOutReconfModuleIRQs_o_0[0]
wire cell_30_0; // PORT

// CellOutReconfModuleIRQs_o_1[0]
wire cell_31_0; // PORT

// CellOutReconfModuleIRQs_o_2[0]
wire cell_32_0; // PORT

// CellOutReconfModuleIRQs_o_3[0]
wire cell_33_0; // PORT

// CellOutReconfModuleIRQs_o_4[0]
wire cell_34_0; // PORT

// CellOutSPI_CPHA_o[0]
wire cell_35_0; // PORT

// CellOutSPI_CPOL_o[0]
wire cell_36_0; // PORT

// CellOutSPI_DataIn_o[0]
wire [7:0] cell_37_0; // PORT

// CellInSPI_DataOut_i[0]
wire [7:0] cell_38_0; // PORT

// CellInSPI_FIFOEmpty_i[0]
wire cell_39_0; // PORT

// CellInSPI_FIFOFull_i[0]
wire cell_40_0; // PORT

// CellOutSPI_LSBFE_o[0]
wire cell_41_0; // PORT

// CellOutSPI_ReadNext_o[0]
wire cell_42_0; // PORT

// CellInSPI_Transmission_i[0]
wire cell_43_0; // PORT

// CellOutSPI_Write_o[0]
wire cell_44_0; // PORT

// CellInReconfModuleIn_i_0[0]
wire cell_45_0; // PORT

// CellInReconfModuleIn_i_1[0]
wire cell_46_0; // PORT

// CellInReconfModuleIn_i_2[0]
wire cell_47_0; // PORT

// CellInReconfModuleIn_i_3[0]
wire cell_48_0; // PORT

// CellInReconfModuleIn_i_4[0]
wire cell_49_0; // PORT

// CellInReconfModuleIn_i_5[0]
wire cell_50_0; // PORT

// CellInReconfModuleIn_i_6[0]
wire cell_51_0; // PORT

// CellInReconfModuleIn_i_7[0]
wire cell_52_0; // PORT

// CellOutReconfModuleOut_o_0[0]
wire cell_53_0; // PORT

// CellOutReconfModuleOut_o_1[0]
wire cell_54_0; // PORT

// CellOutReconfModuleOut_o_2[0]
wire cell_55_0; // PORT

// CellOutReconfModuleOut_o_3[0]
wire cell_56_0; // PORT

// CellOutReconfModuleOut_o_4[0]
wire cell_57_0; // PORT

// CellOutReconfModuleOut_o_5[0]
wire cell_58_0; // PORT

// CellOutReconfModuleOut_o_6[0]
wire cell_59_0; // PORT

// CellOutReconfModuleOut_o_7[0]
wire cell_60_0; // PORT

// Counter[0]
wire [15:0] cell_61_5; // D_o
wire cell_61_3; // Direction_i
wire cell_61_2; // Enable_i
wire cell_61_6; // Overflow_o
wire [15:0] cell_61_4; // PresetVal_i
wire cell_61_1; // Preset_i
wire cell_61_0; // ResetSig_i
wire cell_61_7; // Zero_o
Counter cell_61 (
	.D_o(cell_61_5),
	.Direction_i(cell_61_3),
	.Enable_i(cell_61_2),
	.Overflow_o(cell_61_6),
	.PresetVal_i(cell_61_4),
	.Preset_i(cell_61_1),
	.ResetSig_i(cell_61_0),
	.Zero_o(cell_61_7),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// Counter[1]
wire [15:0] cell_62_5; // D_o
wire cell_62_3; // Direction_i
wire cell_62_2; // Enable_i
wire cell_62_6; // Overflow_o
wire [15:0] cell_62_4; // PresetVal_i
wire cell_62_1; // Preset_i
wire cell_62_0; // ResetSig_i
wire cell_62_7; // Zero_o
Counter cell_62 (
	.D_o(cell_62_5),
	.Direction_i(cell_62_3),
	.Enable_i(cell_62_2),
	.Overflow_o(cell_62_6),
	.PresetVal_i(cell_62_4),
	.Preset_i(cell_62_1),
	.ResetSig_i(cell_62_0),
	.Zero_o(cell_62_7),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// Counter32[0]
wire [15:0] cell_63_6; // DH_o
wire [15:0] cell_63_7; // DL_o
wire cell_63_3; // Direction_i
wire cell_63_2; // Enable_i
wire cell_63_8; // Overflow_o
wire [15:0] cell_63_4; // PresetValH_i
wire [15:0] cell_63_5; // PresetValL_i
wire cell_63_1; // Preset_i
wire cell_63_0; // ResetSig_i
wire cell_63_9; // Zero_o
Counter32 cell_63 (
	.DH_o(cell_63_6),
	.DL_o(cell_63_7),
	.Direction_i(cell_63_3),
	.Enable_i(cell_63_2),
	.Overflow_o(cell_63_8),
	.PresetValH_i(cell_63_4),
	.PresetValL_i(cell_63_5),
	.Preset_i(cell_63_1),
	.ResetSig_i(cell_63_0),
	.Zero_o(cell_63_9),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// Counter32[1]
wire [15:0] cell_64_6; // DH_o
wire [15:0] cell_64_7; // DL_o
wire cell_64_3; // Direction_i
wire cell_64_2; // Enable_i
wire cell_64_8; // Overflow_o
wire [15:0] cell_64_4; // PresetValH_i
wire [15:0] cell_64_5; // PresetValL_i
wire cell_64_1; // Preset_i
wire cell_64_0; // ResetSig_i
wire cell_64_9; // Zero_o
Counter32 cell_64 (
	.DH_o(cell_64_6),
	.DL_o(cell_64_7),
	.Direction_i(cell_64_3),
	.Enable_i(cell_64_2),
	.Overflow_o(cell_64_8),
	.PresetValH_i(cell_64_4),
	.PresetValL_i(cell_64_5),
	.Preset_i(cell_64_1),
	.ResetSig_i(cell_64_0),
	.Zero_o(cell_64_9),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// AbsDiff[0]
wire [15:0] cell_65_0; // A_i
wire [15:0] cell_65_1; // B_i
wire [15:0] cell_65_2; // D_o
AbsDiff cell_65 (
	.A_i(cell_65_0),
	.B_i(cell_65_1),
	.D_o(cell_65_2)
);

// WordRegister[0]
wire [15:0] cell_66_0; // D_i
wire cell_66_2; // Enable_i
wire [15:0] cell_66_1; // Q_o
WordRegister cell_66 (
	.D_i(cell_66_0),
	.Enable_i(cell_66_2),
	.Q_o(cell_66_1),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// WordRegister[1]
wire [15:0] cell_67_0; // D_i
wire cell_67_2; // Enable_i
wire [15:0] cell_67_1; // Q_o
WordRegister cell_67 (
	.D_i(cell_67_0),
	.Enable_i(cell_67_2),
	.Q_o(cell_67_1),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// WordRegister[2]
wire [15:0] cell_68_0; // D_i
wire cell_68_2; // Enable_i
wire [15:0] cell_68_1; // Q_o
WordRegister cell_68 (
	.D_i(cell_68_0),
	.Enable_i(cell_68_2),
	.Q_o(cell_68_1),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// ByteRegister[0]
wire [7:0] cell_69_0; // D_i
wire cell_69_2; // Enable_i
wire [7:0] cell_69_1; // Q_o
ByteRegister cell_69 (
	.D_i(cell_69_0),
	.Enable_i(cell_69_2),
	.Q_o(cell_69_1),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// ByteRegister[1]
wire [7:0] cell_70_0; // D_i
wire cell_70_2; // Enable_i
wire [7:0] cell_70_1; // Q_o
ByteRegister cell_70 (
	.D_i(cell_70_0),
	.Enable_i(cell_70_2),
	.Q_o(cell_70_1),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i)
);

// AddSubCmp[0]
wire [15:0] cell_71_1; // A_i
wire cell_71_0; // AddOrSub_i
wire [15:0] cell_71_2; // B_i
wire cell_71_4; // Carry_i
wire cell_71_5; // Carry_o
wire [15:0] cell_71_3; // D_o
wire cell_71_8; // Overflow_o
wire cell_71_7; // Sign_o
wire cell_71_6; // Zero_o
AddSubCmp cell_71 (
	.A_i(cell_71_1),
	.AddOrSub_i(cell_71_0),
	.B_i(cell_71_2),
	.Carry_i(cell_71_4),
	.Carry_o(cell_71_5),
	.D_o(cell_71_3),
	.Overflow_o(cell_71_8),
	.Sign_o(cell_71_7),
	.Zero_o(cell_71_6)
);

// AddSubCmp[1]
wire [15:0] cell_72_1; // A_i
wire cell_72_0; // AddOrSub_i
wire [15:0] cell_72_2; // B_i
wire cell_72_4; // Carry_i
wire cell_72_5; // Carry_o
wire [15:0] cell_72_3; // D_o
wire cell_72_8; // Overflow_o
wire cell_72_7; // Sign_o
wire cell_72_6; // Zero_o
AddSubCmp cell_72 (
	.A_i(cell_72_1),
	.AddOrSub_i(cell_72_0),
	.B_i(cell_72_2),
	.Carry_i(cell_72_4),
	.Carry_o(cell_72_5),
	.D_o(cell_72_3),
	.Overflow_o(cell_72_8),
	.Sign_o(cell_72_7),
	.Zero_o(cell_72_6)
);

// ByteMuxQuad[0]
wire [7:0] cell_73_0; // A_i
wire [7:0] cell_73_1; // B_i
wire [7:0] cell_73_2; // C_i
wire [7:0] cell_73_3; // D_i
wire cell_73_4; // SAB_i
wire cell_73_5; // SC_i
wire cell_73_6; // SD_i
wire [7:0] cell_73_7; // Y_o
ByteMuxQuad cell_73 (
	.A_i(cell_73_0),
	.B_i(cell_73_1),
	.C_i(cell_73_2),
	.D_i(cell_73_3),
	.SAB_i(cell_73_4),
	.SC_i(cell_73_5),
	.SD_i(cell_73_6),
	.Y_o(cell_73_7)
);

// ByteMuxDual[0]
wire [7:0] cell_74_0; // A_i
wire [7:0] cell_74_1; // B_i
wire cell_74_2; // S_i
wire [7:0] cell_74_3; // Y_o
ByteMuxDual cell_74 (
	.A_i(cell_74_0),
	.B_i(cell_74_1),
	.S_i(cell_74_2),
	.Y_o(cell_74_3)
);

// ByteMuxDual[1]
wire [7:0] cell_75_0; // A_i
wire [7:0] cell_75_1; // B_i
wire cell_75_2; // S_i
wire [7:0] cell_75_3; // Y_o
ByteMuxDual cell_75 (
	.A_i(cell_75_0),
	.B_i(cell_75_1),
	.S_i(cell_75_2),
	.Y_o(cell_75_3)
);

// Byte2Word[0]
wire [7:0] cell_76_0; // H_i
wire [7:0] cell_76_1; // L_i
wire [15:0] cell_76_2; // Y_o
Byte2Word cell_76 (
	.H_i(cell_76_0),
	.L_i(cell_76_1),
	.Y_o(cell_76_2)
);

// Byte2WordSel[0]
wire [7:0] cell_77_0; // H_i
wire [7:0] cell_77_1; // L_i
wire [15:0] cell_77_2; // Y_o
Byte2WordSel cell_77 (
	.H_i(cell_77_0),
	.L_i(cell_77_1),
	.Y_o(cell_77_2),
	.Mask_i(bitdata[1215:1212]),
	.Shift_i(bitdata[1211:1208])
);

// WordMuxDual[0]
wire [15:0] cell_78_0; // A_i
wire [15:0] cell_78_1; // B_i
wire cell_78_2; // S_i
wire [15:0] cell_78_3; // Y_o
WordMuxDual cell_78 (
	.A_i(cell_78_0),
	.B_i(cell_78_1),
	.S_i(cell_78_2),
	.Y_o(cell_78_3)
);

// WordMuxDual[1]
wire [15:0] cell_79_0; // A_i
wire [15:0] cell_79_1; // B_i
wire cell_79_2; // S_i
wire [15:0] cell_79_3; // Y_o
WordMuxDual cell_79 (
	.A_i(cell_79_0),
	.B_i(cell_79_1),
	.S_i(cell_79_2),
	.Y_o(cell_79_3)
);

// TRFSM0[0]
wire cell_80_0; // In0_i
wire cell_80_1; // In1_i
wire cell_80_2; // In2_i
wire cell_80_3; // In3_i
wire cell_80_4; // In4_i
wire cell_80_5; // In5_i
wire cell_80_6; // Out0_o
wire cell_80_7; // Out1_o
wire cell_80_8; // Out2_o
wire cell_80_9; // Out3_o
wire cell_80_10; // Out4_o
wire cell_80_11; // Out5_o
wire cell_80_12; // Out6_o
wire cell_80_13; // Out7_o
wire cell_80_14; // Out8_o
wire cell_80_15; // Out9_o
TRFSM0 cell_80 (
	.In0_i(cell_80_0),
	.In1_i(cell_80_1),
	.In2_i(cell_80_2),
	.In3_i(cell_80_3),
	.In4_i(cell_80_4),
	.In5_i(cell_80_5),
	.Out0_o(cell_80_6),
	.Out1_o(cell_80_7),
	.Out2_o(cell_80_8),
	.Out3_o(cell_80_9),
	.Out4_o(cell_80_10),
	.Out5_o(cell_80_11),
	.Out6_o(cell_80_12),
	.Out7_o(cell_80_13),
	.Out8_o(cell_80_14),
	.Out9_o(cell_80_15),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i),
	.CfgMode_i(CfgMode_i),
	.CfgClk_i(CfgClk_TRFSM0_i),
	.CfgShift_i(CfgShift_TRFSM0_i),
	.CfgDataIn_i(CfgDataIn_i),
	.CfgDataOut_o(CfgDataOut_TRFSM0_o)
);

// TRFSM1[0]
wire cell_81_0; // In0_i
wire cell_81_1; // In1_i
wire cell_81_2; // In2_i
wire cell_81_3; // In3_i
wire cell_81_4; // In4_i
wire cell_81_5; // In5_i
wire cell_81_6; // In6_i
wire cell_81_7; // In7_i
wire cell_81_8; // In8_i
wire cell_81_9; // In9_i
wire cell_81_10; // Out0_o
wire cell_81_20; // Out10_o
wire cell_81_21; // Out11_o
wire cell_81_22; // Out12_o
wire cell_81_23; // Out13_o
wire cell_81_24; // Out14_o
wire cell_81_11; // Out1_o
wire cell_81_12; // Out2_o
wire cell_81_13; // Out3_o
wire cell_81_14; // Out4_o
wire cell_81_15; // Out5_o
wire cell_81_16; // Out6_o
wire cell_81_17; // Out7_o
wire cell_81_18; // Out8_o
wire cell_81_19; // Out9_o
TRFSM1 cell_81 (
	.In0_i(cell_81_0),
	.In1_i(cell_81_1),
	.In2_i(cell_81_2),
	.In3_i(cell_81_3),
	.In4_i(cell_81_4),
	.In5_i(cell_81_5),
	.In6_i(cell_81_6),
	.In7_i(cell_81_7),
	.In8_i(cell_81_8),
	.In9_i(cell_81_9),
	.Out0_o(cell_81_10),
	.Out10_o(cell_81_20),
	.Out11_o(cell_81_21),
	.Out12_o(cell_81_22),
	.Out13_o(cell_81_23),
	.Out14_o(cell_81_24),
	.Out1_o(cell_81_11),
	.Out2_o(cell_81_12),
	.Out3_o(cell_81_13),
	.Out4_o(cell_81_14),
	.Out5_o(cell_81_15),
	.Out6_o(cell_81_16),
	.Out7_o(cell_81_17),
	.Out8_o(cell_81_18),
	.Out9_o(cell_81_19),
	.Clk_i(Clk_i),
	.Reset_n_i(Reset_n_i),
	.CfgMode_i(CfgMode_i),
	.CfgClk_i(CfgClk_TRFSM1_i),
	.CfgShift_i(CfgShift_TRFSM1_i),
	.CfgDataIn_i(CfgDataIn_i),
	.CfgDataOut_o(CfgDataOut_TRFSM1_o)
);

// CONST_Bit[0]
wire cell_82_0; // Value_o
CONST_Bit cell_82 (
	.Value_o(cell_82_0),
	.CfgValue_i(bitdata[1216:1216])
);

// CONST_Bit[1]
wire cell_83_0; // Value_o
CONST_Bit cell_83 (
	.Value_o(cell_83_0),
	.CfgValue_i(bitdata[1217:1217])
);

// CONST_Byte[0]
wire [7:0] cell_84_0; // Value_o
CONST_Byte cell_84 (
	.Value_o(cell_84_0),
	.CfgValue_i(bitdata[1225:1218])
);

// CONST_Byte[1]
wire [7:0] cell_85_0; // Value_o
CONST_Byte cell_85 (
	.Value_o(cell_85_0),
	.CfgValue_i(bitdata[1233:1226])
);

// CONST_Byte[2]
wire [7:0] cell_86_0; // Value_o
CONST_Byte cell_86 (
	.Value_o(cell_86_0),
	.CfgValue_i(bitdata[1241:1234])
);

// CONST_Byte[3]
wire [7:0] cell_87_0; // Value_o
CONST_Byte cell_87 (
	.Value_o(cell_87_0),
	.CfgValue_i(bitdata[1249:1242])
);

// CONST_Byte[4]
wire [7:0] cell_88_0; // Value_o
CONST_Byte cell_88 (
	.Value_o(cell_88_0),
	.CfgValue_i(bitdata[1257:1250])
);

// CONST_Byte[5]
wire [7:0] cell_89_0; // Value_o
CONST_Byte cell_89 (
	.Value_o(cell_89_0),
	.CfgValue_i(bitdata[1265:1258])
);

// CONST_Word[0]
wire [15:0] cell_90_0; // Value_o
CONST_Word cell_90 (
	.Value_o(cell_90_0),
	.CfgValue_i(bitdata[1281:1266])
);

// CellParamIn_Word[0]
wire [15:0] cell_91_0; // PORT

// CellParamIn_Word[1]
wire [15:0] cell_92_0; // PORT

// CellParamIn_Word[2]
wire [15:0] cell_93_0; // PORT

// CellParamIn_Word[3]
wire [15:0] cell_94_0; // PORT

// CellParamIn_Word[4]
wire [15:0] cell_95_0; // PORT

// CellParamOut_Word[0]
wire [15:0] cell_96_0; // PORT

// CellParamOut_Word[1]
wire [15:0] cell_97_0; // PORT

// input and output mappings to interconnect signals
assign cell_0_0 = AdcConvComplete_i;
assign AdcDoConvert_o = cell_1_0;
assign cell_2_0 = AdcValue_i;
assign cell_3_0 = I2C_Busy_i;
assign I2C_DataIn_o = cell_4_0;
assign cell_5_0 = I2C_DataOut_i;
assign cell_6_0 = I2C_Error_i;
assign cell_7_0 = I2C_FIFOEmpty_i;
assign cell_8_0 = I2C_FIFOFull_i;
assign I2C_FIFOReadNext_o = cell_9_0;
assign I2C_FIFOWrite_o = cell_10_0;
assign I2C_ReadCount_o = cell_11_0;
assign I2C_ReceiveSend_n_o = cell_12_0;
assign I2C_StartProcess_o = cell_13_0;
assign cell_14_0 = Inputs_i_0;
assign cell_15_0 = Inputs_i_1;
assign cell_16_0 = Inputs_i_2;
assign cell_17_0 = Inputs_i_3;
assign cell_18_0 = Inputs_i_4;
assign cell_19_0 = Inputs_i_5;
assign cell_20_0 = Inputs_i_6;
assign cell_21_0 = Inputs_i_7;
assign Outputs_o_0 = cell_22_0;
assign Outputs_o_1 = cell_23_0;
assign Outputs_o_2 = cell_24_0;
assign Outputs_o_3 = cell_25_0;
assign Outputs_o_4 = cell_26_0;
assign Outputs_o_5 = cell_27_0;
assign Outputs_o_6 = cell_28_0;
assign Outputs_o_7 = cell_29_0;
assign ReconfModuleIRQs_o_0 = cell_30_0;
assign ReconfModuleIRQs_o_1 = cell_31_0;
assign ReconfModuleIRQs_o_2 = cell_32_0;
assign ReconfModuleIRQs_o_3 = cell_33_0;
assign ReconfModuleIRQs_o_4 = cell_34_0;
assign SPI_CPHA_o = cell_35_0;
assign SPI_CPOL_o = cell_36_0;
assign SPI_DataIn_o = cell_37_0;
assign cell_38_0 = SPI_DataOut_i;
assign cell_39_0 = SPI_FIFOEmpty_i;
assign cell_40_0 = SPI_FIFOFull_i;
assign SPI_LSBFE_o = cell_41_0;
assign SPI_ReadNext_o = cell_42_0;
assign cell_43_0 = SPI_Transmission_i;
assign SPI_Write_o = cell_44_0;
assign cell_45_0 = ReconfModuleIn_i_0;
assign cell_46_0 = ReconfModuleIn_i_1;
assign cell_47_0 = ReconfModuleIn_i_2;
assign cell_48_0 = ReconfModuleIn_i_3;
assign cell_49_0 = ReconfModuleIn_i_4;
assign cell_50_0 = ReconfModuleIn_i_5;
assign cell_51_0 = ReconfModuleIn_i_6;
assign cell_52_0 = ReconfModuleIn_i_7;
assign ReconfModuleOut_o_0 = cell_53_0;
assign ReconfModuleOut_o_1 = cell_54_0;
assign ReconfModuleOut_o_2 = cell_55_0;
assign ReconfModuleOut_o_3 = cell_56_0;
assign ReconfModuleOut_o_4 = cell_57_0;
assign ReconfModuleOut_o_5 = cell_58_0;
assign ReconfModuleOut_o_6 = cell_59_0;
assign ReconfModuleOut_o_7 = cell_60_0;
assign cell_91_0 = ParamIn_Word_i[15:0];
assign cell_92_0 = ParamIn_Word_i[31:16];
assign cell_93_0 = ParamIn_Word_i[47:32];
assign cell_94_0 = ParamIn_Word_i[63:48];
assign cell_95_0 = ParamIn_Word_i[79:64];
assign ParamOut_Word_o[15:0] = cell_96_0;
assign ParamOut_Word_o[31:16] = cell_97_0;

// conntype=0, tree=0, switch=1
wire sw_0_0_1_up0;
wire sw_0_0_1_down0;

// conntype=0, tree=0, switch=2
wire sw_0_0_2_up0;
wire sw_0_0_2_down0;

// conntype=0, tree=0, switch=3
wire sw_0_0_3_up0;
wire sw_0_0_3_down0;

// conntype=0, tree=0, switch=4
wire sw_0_0_4_up0;
wire sw_0_0_4_down0;

// conntype=0, tree=0, switch=5
wire sw_0_0_5_up0;
wire sw_0_0_5_down0;

// conntype=0, tree=0, switch=6
wire sw_0_0_6_up0;
wire sw_0_0_6_down0;

// conntype=0, tree=0, switch=7
wire sw_0_0_7_up0;
wire sw_0_0_7_down0;

// conntype=0, tree=0, switch=8
wire sw_0_0_8_up0;
wire sw_0_0_8_up1;
wire sw_0_0_8_up2;
wire sw_0_0_8_down0;
wire sw_0_0_8_down1;
wire sw_0_0_8_down2;
wire sw_0_0_8_down3;
wire sw_0_0_8_down4;

// conntype=0, tree=0, switch=9
wire sw_0_0_9_up0;
wire sw_0_0_9_up1;
wire sw_0_0_9_up2;
wire sw_0_0_9_up3;

// conntype=0, tree=0, switch=10
wire sw_0_0_10_up0;
wire sw_0_0_10_down0;
wire sw_0_0_10_down1;
wire sw_0_0_10_down2;

// conntype=0, tree=0, switch=11
wire sw_0_0_11_up0;
wire sw_0_0_11_down0;
wire sw_0_0_11_down1;

// conntype=0, tree=0, switch=12
wire sw_0_0_12_up0;
wire sw_0_0_12_down0;

// conntype=0, tree=0, switch=13
wire sw_0_0_13_down0;

// conntype=0, tree=0, switch=14
wire sw_0_0_14_down0;

// conntype=0, tree=0, switch=15
wire sw_0_0_15_up0;

// conntype=0, tree=0, switch=16
wire sw_0_0_16_up0;
wire sw_0_0_16_down0;

// conntype=0, tree=0, switch=17
wire sw_0_0_17_down0;

// conntype=0, tree=0, switch=18
wire sw_0_0_18_up0;
wire sw_0_0_18_down0;

// conntype=0, tree=0, switch=19
wire sw_0_0_19_down0;

// conntype=0, tree=0, switch=20
wire sw_0_0_20_up0;
wire sw_0_0_20_down0;

// conntype=0, tree=0, switch=21
wire sw_0_0_21_down0;

// conntype=0, tree=0, switch=22
wire sw_0_0_22_up0;
wire sw_0_0_22_down0;

// conntype=0, tree=0, switch=23
wire sw_0_0_23_up0;

// conntype=0, tree=0, switch=24
wire sw_0_0_24_up0;
wire sw_0_0_24_down0;
wire sw_0_0_24_down1;
wire sw_0_0_24_down2;

// conntype=0, tree=0, switch=25
wire sw_0_0_25_up0;
wire sw_0_0_25_up1;
wire sw_0_0_25_up2;
wire sw_0_0_25_up3;
wire sw_0_0_25_down0;
wire sw_0_0_25_down1;
wire sw_0_0_25_down2;

// conntype=0, tree=0, switch=26
wire sw_0_0_26_up0;
wire sw_0_0_26_down0;
wire sw_0_0_26_down1;

// conntype=0, tree=1, switch=1
wire sw_0_1_1_up0;
wire sw_0_1_1_down0;

// conntype=0, tree=1, switch=2
wire sw_0_1_2_up0;
wire sw_0_1_2_down0;

// conntype=0, tree=1, switch=3
wire sw_0_1_3_up0;
wire sw_0_1_3_up1;
wire sw_0_1_3_up2;
wire sw_0_1_3_up3;
wire sw_0_1_3_up4;
wire sw_0_1_3_up5;
wire sw_0_1_3_down0;
wire sw_0_1_3_down1;

// conntype=0, tree=1, switch=4
wire sw_0_1_4_up0;
wire sw_0_1_4_down0;
wire sw_0_1_4_down1;

// conntype=0, tree=1, switch=5
wire sw_0_1_5_up0;
wire sw_0_1_5_up1;
wire sw_0_1_5_down0;
wire sw_0_1_5_down1;
wire sw_0_1_5_down2;
wire sw_0_1_5_down3;
wire sw_0_1_5_down4;

// conntype=0, tree=1, switch=6
wire sw_0_1_6_up0;
wire sw_0_1_6_down0;

// conntype=0, tree=1, switch=7
wire sw_0_1_7_up0;
wire sw_0_1_7_down0;

// conntype=0, tree=1, switch=8
wire sw_0_1_8_up0;
wire sw_0_1_8_up1;
wire sw_0_1_8_up2;
wire sw_0_1_8_up3;
wire sw_0_1_8_up4;
wire sw_0_1_8_up5;
wire sw_0_1_8_up6;
wire sw_0_1_8_up7;
wire sw_0_1_8_up8;
wire sw_0_1_8_up9;
wire sw_0_1_8_down0;
wire sw_0_1_8_down1;
wire sw_0_1_8_down2;
wire sw_0_1_8_down3;
wire sw_0_1_8_down4;
wire sw_0_1_8_down5;

// conntype=0, tree=1, switch=9
wire sw_0_1_9_up0;
wire sw_0_1_9_down0;
wire sw_0_1_9_down1;
wire sw_0_1_9_down2;

// conntype=0, tree=1, switch=10
wire sw_0_1_10_up0;
wire sw_0_1_10_up1;
wire sw_0_1_10_up2;
wire sw_0_1_10_down0;
wire sw_0_1_10_down1;
wire sw_0_1_10_down2;
wire sw_0_1_10_down3;
wire sw_0_1_10_down4;

// conntype=0, tree=1, switch=11
wire sw_0_1_11_up0;
wire sw_0_1_11_up1;
wire sw_0_1_11_up2;
wire sw_0_1_11_up3;
wire sw_0_1_11_down0;
wire sw_0_1_11_down1;
wire sw_0_1_11_down2;
wire sw_0_1_11_down3;

// conntype=0, tree=1, switch=12
wire sw_0_1_12_down0;
wire sw_0_1_12_down1;

// conntype=0, tree=1, switch=13
wire sw_0_1_13_down0;

// conntype=0, tree=1, switch=14
wire sw_0_1_14_down0;

// conntype=0, tree=1, switch=15
wire sw_0_1_15_up0;

// conntype=0, tree=1, switch=16
wire sw_0_1_16_up0;
wire sw_0_1_16_up1;

// conntype=0, tree=1, switch=17
wire sw_0_1_17_up0;
wire sw_0_1_17_down0;
wire sw_0_1_17_down1;
wire sw_0_1_17_down2;

// conntype=0, tree=1, switch=18
wire sw_0_1_18_up0;
wire sw_0_1_18_down0;
wire sw_0_1_18_down1;
wire sw_0_1_18_down2;

// conntype=0, tree=1, switch=19
wire sw_0_1_19_up0;
wire sw_0_1_19_down0;
wire sw_0_1_19_down1;

// conntype=0, tree=1, switch=20
wire sw_0_1_20_down0;

// conntype=0, tree=1, switch=21
wire sw_0_1_21_down0;

// conntype=0, tree=1, switch=22
wire sw_0_1_22_up0;
wire sw_0_1_22_down0;

// conntype=0, tree=1, switch=23
wire sw_0_1_23_up0;

// conntype=0, tree=1, switch=24
wire sw_0_1_24_up0;
wire sw_0_1_24_down0;

// conntype=0, tree=1, switch=25
wire sw_0_1_25_up0;
wire sw_0_1_25_down0;

// conntype=0, tree=1, switch=26
wire sw_0_1_26_up0;
wire sw_0_1_26_down0;

// conntype=1, tree=0, switch=1
wire [7:0] sw_1_0_1_up0;
wire [7:0] sw_1_0_1_down0;

// conntype=1, tree=0, switch=2
wire [7:0] sw_1_0_2_up0;
wire [7:0] sw_1_0_2_down0;

// conntype=1, tree=0, switch=3
wire [7:0] sw_1_0_3_up0;
wire [7:0] sw_1_0_3_down0;
wire [7:0] sw_1_0_3_down1;

// conntype=1, tree=0, switch=4
wire [7:0] sw_1_0_4_up0;
wire [7:0] sw_1_0_4_up1;
wire [7:0] sw_1_0_4_down0;

// conntype=1, tree=0, switch=5
wire [7:0] sw_1_0_5_up0;
wire [7:0] sw_1_0_5_down0;

// conntype=1, tree=0, switch=6
wire [7:0] sw_1_0_6_up0;
wire [7:0] sw_1_0_6_down0;

// conntype=1, tree=0, switch=7
wire [7:0] sw_1_0_7_up0;

// conntype=1, tree=1, switch=1
wire [7:0] sw_1_1_1_up0;
wire [7:0] sw_1_1_1_down0;

// conntype=1, tree=1, switch=2
wire [7:0] sw_1_1_2_up0;
wire [7:0] sw_1_1_2_down0;

// conntype=1, tree=1, switch=3
wire [7:0] sw_1_1_3_up0;
wire [7:0] sw_1_1_3_down0;

// conntype=1, tree=1, switch=4
wire [7:0] sw_1_1_4_up0;
wire [7:0] sw_1_1_4_up1;
wire [7:0] sw_1_1_4_down0;

// conntype=1, tree=1, switch=5
wire [7:0] sw_1_1_5_up0;
wire [7:0] sw_1_1_5_down0;
wire [7:0] sw_1_1_5_down1;

// conntype=1, tree=1, switch=6
wire [7:0] sw_1_1_6_up0;
wire [7:0] sw_1_1_6_down0;

// conntype=1, tree=1, switch=7
wire [7:0] sw_1_1_7_down0;

// conntype=2, tree=0, switch=1
wire [15:0] sw_2_0_1_up0;
wire [15:0] sw_2_0_1_down0;

// conntype=2, tree=0, switch=2
wire [15:0] sw_2_0_2_up0;
wire [15:0] sw_2_0_2_down0;

// conntype=2, tree=0, switch=3
wire [15:0] sw_2_0_3_up0;
wire [15:0] sw_2_0_3_down0;

// conntype=2, tree=0, switch=4
wire [15:0] sw_2_0_4_up0;
wire [15:0] sw_2_0_4_down0;

// conntype=2, tree=0, switch=5
wire [15:0] sw_2_0_5_up0;
wire [15:0] sw_2_0_5_down0;

// conntype=2, tree=0, switch=6
wire [15:0] sw_2_0_6_up0;
wire [15:0] sw_2_0_6_down0;

// conntype=2, tree=0, switch=7
wire [15:0] sw_2_0_7_up0;
wire [15:0] sw_2_0_7_down0;

// conntype=2, tree=0, switch=8
wire [15:0] sw_2_0_8_up0;
wire [15:0] sw_2_0_8_down0;

// conntype=2, tree=1, switch=1
wire [15:0] sw_2_1_1_up0;
wire [15:0] sw_2_1_1_down0;

// conntype=2, tree=1, switch=2
wire [15:0] sw_2_1_2_up0;
wire [15:0] sw_2_1_2_down0;

// conntype=2, tree=1, switch=3
wire [15:0] sw_2_1_3_up0;
wire [15:0] sw_2_1_3_down0;

// conntype=2, tree=1, switch=4
wire [15:0] sw_2_1_4_up0;
wire [15:0] sw_2_1_4_down0;

// conntype=2, tree=1, switch=5
wire [15:0] sw_2_1_5_up0;
wire [15:0] sw_2_1_5_down0;

// conntype=2, tree=1, switch=6
wire [15:0] sw_2_1_6_up0;
wire [15:0] sw_2_1_6_up1;
wire [15:0] sw_2_1_6_down0;

// conntype=2, tree=1, switch=7
wire [15:0] sw_2_1_7_up0;
wire [15:0] sw_2_1_7_down0;
wire [15:0] sw_2_1_7_down1;

// conntype=2, tree=1, switch=8
wire [15:0] sw_2_1_8_up0;
wire [15:0] sw_2_1_8_down0;

// multiplexer
assign cell_10_0 =
   (bitdata[271:269] == 3'b010 ? sw_0_0_24_down0 :
    bitdata[271:269] == 3'b110 ? sw_0_0_24_down1 :
    bitdata[271:269] == 3'b001 ? sw_0_0_24_down2 :
    bitdata[271:269] == 3'b100 ? cell_3_0 :
    bitdata[271:269] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[898:897] == 2'b01 ? sw_0_1_24_down0 :
    bitdata[898:897] == 2'b10 ? cell_14_0 :
    bitdata[898:897] == 2'b0 ? 1'b0 : 1'bx);
assign cell_11_0 =
   (bitdata[946:944] == 3'b001 ? sw_1_0_4_down0 :
    bitdata[946:944] == 3'b100 ? cell_74_3 :
    bitdata[946:944] == 3'b010 ? cell_84_0 :
    bitdata[946:944] == 3'b110 ? cell_85_0 :
    bitdata[946:944] == 3'b0 ? 8'b0 : 8'bx) |
   (bitdata[1031:1031] == 1'b1 ? sw_1_1_7_down0 :
    bitdata[1031:1031] == 1'b0 ? 8'b0 : 8'bx);
assign cell_12_0 =
   (bitdata[369:368] == 2'b01 ? sw_0_0_26_down0 :
    bitdata[369:368] == 2'b11 ? sw_0_0_26_down1 :
    bitdata[369:368] == 2'b10 ? cell_6_0 :
    bitdata[369:368] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[900:899] == 2'b01 ? sw_0_1_24_down0 :
    bitdata[900:899] == 2'b10 ? cell_14_0 :
    bitdata[900:899] == 2'b0 ? 1'b0 : 1'bx);
assign cell_13_0 =
   (bitdata[274:272] == 3'b010 ? sw_0_0_24_down0 :
    bitdata[274:272] == 3'b110 ? sw_0_0_24_down1 :
    bitdata[274:272] == 3'b001 ? sw_0_0_24_down2 :
    bitdata[274:272] == 3'b100 ? cell_3_0 :
    bitdata[274:272] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[902:901] == 2'b01 ? sw_0_1_24_down0 :
    bitdata[902:901] == 2'b10 ? cell_14_0 :
    bitdata[902:901] == 2'b0 ? 1'b0 : 1'bx);
assign cell_1_0 =
   (bitdata[180:177] == 4'b0110 ? sw_0_0_10_down0 :
    bitdata[180:177] == 4'b1110 ? sw_0_0_10_down1 :
    bitdata[180:177] == 4'b0001 ? sw_0_0_10_down2 :
    bitdata[180:177] == 4'b1000 ? cell_62_6 :
    bitdata[180:177] == 4'b0100 ? cell_62_7 :
    bitdata[180:177] == 4'b1100 ? cell_64_8 :
    bitdata[180:177] == 4'b0010 ? cell_64_9 :
    bitdata[180:177] == 4'b1010 ? cell_83_0 :
    bitdata[180:177] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[910:909] == 2'b11 ? sw_0_1_26_down0 :
    bitdata[910:909] == 2'b10 ? cell_0_0 :
    bitdata[910:909] == 2'b01 ? cell_3_0 :
    bitdata[910:909] == 2'b0 ? 1'b0 : 1'bx);
assign cell_22_0 =
   (bitdata[206:205] == 2'b01 ? sw_0_0_11_down0 :
    bitdata[206:205] == 2'b11 ? sw_0_0_11_down1 :
    bitdata[206:205] == 2'b10 ? cell_43_0 :
    bitdata[206:205] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[718:716] == 3'b010 ? sw_0_1_9_down0 :
    bitdata[718:716] == 3'b110 ? sw_0_1_9_down1 :
    bitdata[718:716] == 3'b001 ? sw_0_1_9_down2 :
    bitdata[718:716] == 3'b100 ? cell_43_0 :
    bitdata[718:716] == 3'b0 ? 1'b0 : 1'bx);
assign cell_23_0 =
   (bitdata[208:207] == 2'b01 ? sw_0_0_11_down0 :
    bitdata[208:207] == 2'b11 ? sw_0_0_11_down1 :
    bitdata[208:207] == 2'b10 ? cell_43_0 :
    bitdata[208:207] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[886:886] == 1'b1 ? sw_0_1_21_down0 :
    bitdata[886:886] == 1'b0 ? 1'b0 : 1'bx);
assign cell_24_0 =
   (bitdata[258:258] == 1'b1 ? sw_0_0_21_down0 :
    bitdata[258:258] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[887:887] == 1'b1 ? sw_0_1_21_down0 :
    bitdata[887:887] == 1'b0 ? 1'b0 : 1'bx);
assign cell_25_0 =
   (bitdata[259:259] == 1'b1 ? sw_0_0_21_down0 :
    bitdata[259:259] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[888:888] == 1'b1 ? sw_0_1_21_down0 :
    bitdata[888:888] == 1'b0 ? 1'b0 : 1'bx);
assign cell_26_0 =
   (bitdata[260:260] == 1'b1 ? sw_0_0_21_down0 :
    bitdata[260:260] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[889:889] == 1'b1 ? sw_0_1_21_down0 :
    bitdata[889:889] == 1'b0 ? 1'b0 : 1'bx);
assign cell_27_0 =
   (bitdata[253:252] == 2'b01 ? sw_0_0_20_down0 :
    bitdata[253:252] == 2'b10 ? cell_7_0 :
    bitdata[253:252] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[882:882] == 1'b1 ? sw_0_1_20_down0 :
    bitdata[882:882] == 1'b0 ? 1'b0 : 1'bx);
assign cell_28_0 =
   (bitdata[255:254] == 2'b01 ? sw_0_0_20_down0 :
    bitdata[255:254] == 2'b10 ? cell_7_0 :
    bitdata[255:254] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[883:883] == 1'b1 ? sw_0_1_20_down0 :
    bitdata[883:883] == 1'b0 ? 1'b0 : 1'bx);
assign cell_29_0 =
   (bitdata[257:256] == 2'b01 ? sw_0_0_20_down0 :
    bitdata[257:256] == 2'b10 ? cell_7_0 :
    bitdata[257:256] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[884:884] == 1'b1 ? sw_0_1_20_down0 :
    bitdata[884:884] == 1'b0 ? 1'b0 : 1'bx);
assign cell_30_0 =
   (bitdata[111:107] == 5'b10001 ? sw_0_0_8_down0 :
    bitdata[111:107] == 5'b01001 ? sw_0_0_8_down1 :
    bitdata[111:107] == 5'b11001 ? sw_0_0_8_down2 :
    bitdata[111:107] == 5'b00101 ? sw_0_0_8_down3 :
    bitdata[111:107] == 5'b10101 ? sw_0_0_8_down4 :
    bitdata[111:107] == 5'b10000 ? cell_61_6 :
    bitdata[111:107] == 5'b01000 ? cell_61_7 :
    bitdata[111:107] == 5'b11000 ? cell_71_5 :
    bitdata[111:107] == 5'b00100 ? cell_71_6 :
    bitdata[111:107] == 5'b10100 ? cell_71_7 :
    bitdata[111:107] == 5'b01100 ? cell_71_8 :
    bitdata[111:107] == 5'b11100 ? cell_80_6 :
    bitdata[111:107] == 5'b00010 ? cell_80_7 :
    bitdata[111:107] == 5'b10010 ? cell_80_8 :
    bitdata[111:107] == 5'b01010 ? cell_80_9 :
    bitdata[111:107] == 5'b11010 ? cell_80_10 :
    bitdata[111:107] == 5'b00110 ? cell_80_11 :
    bitdata[111:107] == 5'b10110 ? cell_80_12 :
    bitdata[111:107] == 5'b01110 ? cell_80_13 :
    bitdata[111:107] == 5'b11110 ? cell_80_14 :
    bitdata[111:107] == 5'b00001 ? cell_80_15 :
    bitdata[111:107] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[877:876] == 2'b01 ? sw_0_1_19_down0 :
    bitdata[877:876] == 2'b11 ? sw_0_1_19_down1 :
    bitdata[877:876] == 2'b10 ? cell_40_0 :
    bitdata[877:876] == 2'b0 ? 1'b0 : 1'bx);
assign cell_31_0 =
   (bitdata[248:248] == 1'b1 ? sw_0_0_19_down0 :
    bitdata[248:248] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[894:892] == 3'b001 ? sw_0_1_22_down0 :
    bitdata[894:892] == 3'b100 ? cell_19_0 :
    bitdata[894:892] == 3'b010 ? cell_20_0 :
    bitdata[894:892] == 3'b110 ? cell_21_0 :
    bitdata[894:892] == 3'b0 ? 1'b0 : 1'bx);
assign cell_32_0 =
   (bitdata[249:249] == 1'b1 ? sw_0_0_19_down0 :
    bitdata[249:249] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[885:885] == 1'b1 ? sw_0_1_20_down0 :
    bitdata[885:885] == 1'b0 ? 1'b0 : 1'bx);
assign cell_33_0 =
   (bitdata[250:250] == 1'b1 ? sw_0_0_19_down0 :
    bitdata[250:250] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[879:878] == 2'b01 ? sw_0_1_19_down0 :
    bitdata[879:878] == 2'b11 ? sw_0_1_19_down1 :
    bitdata[879:878] == 2'b10 ? cell_40_0 :
    bitdata[879:878] == 2'b0 ? 1'b0 : 1'bx);
assign cell_34_0 =
   (bitdata[251:251] == 1'b1 ? sw_0_0_19_down0 :
    bitdata[251:251] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[881:880] == 2'b01 ? sw_0_1_19_down0 :
    bitdata[881:880] == 2'b11 ? sw_0_1_19_down1 :
    bitdata[881:880] == 2'b10 ? cell_40_0 :
    bitdata[881:880] == 2'b0 ? 1'b0 : 1'bx);
assign cell_35_0 =
   (bitdata[245:244] == 2'b11 ? sw_0_0_18_down0 :
    bitdata[245:244] == 2'b10 ? cell_39_0 :
    bitdata[245:244] == 2'b01 ? cell_40_0 :
    bitdata[245:244] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[865:863] == 3'b101 ? sw_0_1_18_down0 :
    bitdata[865:863] == 3'b011 ? sw_0_1_18_down1 :
    bitdata[865:863] == 3'b111 ? sw_0_1_18_down2 :
    bitdata[865:863] == 3'b100 ? cell_72_5 :
    bitdata[865:863] == 3'b010 ? cell_72_6 :
    bitdata[865:863] == 3'b110 ? cell_72_7 :
    bitdata[865:863] == 3'b001 ? cell_72_8 :
    bitdata[865:863] == 3'b0 ? 1'b0 : 1'bx);
assign cell_36_0 =
   (bitdata[247:246] == 2'b11 ? sw_0_0_18_down0 :
    bitdata[247:246] == 2'b10 ? cell_39_0 :
    bitdata[247:246] == 2'b01 ? cell_40_0 :
    bitdata[247:246] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[868:866] == 3'b101 ? sw_0_1_18_down0 :
    bitdata[868:866] == 3'b011 ? sw_0_1_18_down1 :
    bitdata[868:866] == 3'b111 ? sw_0_1_18_down2 :
    bitdata[868:866] == 3'b100 ? cell_72_5 :
    bitdata[868:866] == 3'b010 ? cell_72_6 :
    bitdata[868:866] == 3'b110 ? cell_72_7 :
    bitdata[868:866] == 3'b001 ? cell_72_8 :
    bitdata[868:866] == 3'b0 ? 1'b0 : 1'bx);
assign cell_37_0 =
   (bitdata[927:925] == 3'b001 ? sw_1_0_3_down0 :
    bitdata[927:925] == 3'b101 ? sw_1_0_3_down1 :
    bitdata[927:925] == 3'b100 ? cell_73_7 :
    bitdata[927:925] == 3'b010 ? cell_87_0 :
    bitdata[927:925] == 3'b110 ? cell_89_0 :
    bitdata[927:925] == 3'b0 ? 8'b0 : 8'bx) |
   (bitdata[1032:1032] == 1'b1 ? sw_1_1_7_down0 :
    bitdata[1032:1032] == 1'b0 ? 8'b0 : 8'bx);
assign cell_41_0 =
   (bitdata[239:239] == 1'b1 ? sw_0_0_17_down0 :
    bitdata[239:239] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[871:869] == 3'b101 ? sw_0_1_18_down0 :
    bitdata[871:869] == 3'b011 ? sw_0_1_18_down1 :
    bitdata[871:869] == 3'b111 ? sw_0_1_18_down2 :
    bitdata[871:869] == 3'b100 ? cell_72_5 :
    bitdata[871:869] == 3'b010 ? cell_72_6 :
    bitdata[871:869] == 3'b110 ? cell_72_7 :
    bitdata[871:869] == 3'b001 ? cell_72_8 :
    bitdata[871:869] == 3'b0 ? 1'b0 : 1'bx);
assign cell_42_0 =
   (bitdata[277:275] == 3'b010 ? sw_0_0_24_down0 :
    bitdata[277:275] == 3'b110 ? sw_0_0_24_down1 :
    bitdata[277:275] == 3'b001 ? sw_0_0_24_down2 :
    bitdata[277:275] == 3'b100 ? cell_3_0 :
    bitdata[277:275] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[854:852] == 3'b010 ? sw_0_1_17_down0 :
    bitdata[854:852] == 3'b110 ? sw_0_1_17_down1 :
    bitdata[854:852] == 3'b001 ? sw_0_1_17_down2 :
    bitdata[854:852] == 3'b100 ? cell_39_0 :
    bitdata[854:852] == 3'b0 ? 1'b0 : 1'bx);
assign cell_44_0 =
   (bitdata[210:209] == 2'b01 ? sw_0_0_11_down0 :
    bitdata[210:209] == 2'b11 ? sw_0_0_11_down1 :
    bitdata[210:209] == 2'b10 ? cell_43_0 :
    bitdata[210:209] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[721:719] == 3'b010 ? sw_0_1_9_down0 :
    bitdata[721:719] == 3'b110 ? sw_0_1_9_down1 :
    bitdata[721:719] == 3'b001 ? sw_0_1_9_down2 :
    bitdata[721:719] == 3'b100 ? cell_43_0 :
    bitdata[721:719] == 3'b0 ? 1'b0 : 1'bx);
assign cell_4_0 =
   (bitdata[953:952] == 2'b11 ? sw_1_0_5_down0 :
    bitdata[953:952] == 2'b10 ? cell_75_3 :
    bitdata[953:952] == 2'b01 ? cell_86_0 :
    bitdata[953:952] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[1030:1030] == 1'b1 ? sw_1_1_7_down0 :
    bitdata[1030:1030] == 1'b0 ? 8'b0 : 8'bx);
assign cell_53_0 =
   (bitdata[228:228] == 1'b1 ? sw_0_0_14_down0 :
    bitdata[228:228] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[842:842] == 1'b1 ? sw_0_1_14_down0 :
    bitdata[842:842] == 1'b0 ? 1'b0 : 1'bx);
assign cell_54_0 =
   (bitdata[229:229] == 1'b1 ? sw_0_0_14_down0 :
    bitdata[229:229] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[843:843] == 1'b1 ? sw_0_1_14_down0 :
    bitdata[843:843] == 1'b0 ? 1'b0 : 1'bx);
assign cell_55_0 =
   (bitdata[230:230] == 1'b1 ? sw_0_0_14_down0 :
    bitdata[230:230] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[844:844] == 1'b1 ? sw_0_1_14_down0 :
    bitdata[844:844] == 1'b0 ? 1'b0 : 1'bx);
assign cell_56_0 =
   (bitdata[231:231] == 1'b1 ? sw_0_0_14_down0 :
    bitdata[231:231] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[845:845] == 1'b1 ? sw_0_1_14_down0 :
    bitdata[845:845] == 1'b0 ? 1'b0 : 1'bx);
assign cell_57_0 =
   (bitdata[224:224] == 1'b1 ? sw_0_0_13_down0 :
    bitdata[224:224] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[838:838] == 1'b1 ? sw_0_1_13_down0 :
    bitdata[838:838] == 1'b0 ? 1'b0 : 1'bx);
assign cell_58_0 =
   (bitdata[225:225] == 1'b1 ? sw_0_0_13_down0 :
    bitdata[225:225] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[839:839] == 1'b1 ? sw_0_1_13_down0 :
    bitdata[839:839] == 1'b0 ? 1'b0 : 1'bx);
assign cell_59_0 =
   (bitdata[226:226] == 1'b1 ? sw_0_0_13_down0 :
    bitdata[226:226] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[840:840] == 1'b1 ? sw_0_1_13_down0 :
    bitdata[840:840] == 1'b0 ? 1'b0 : 1'bx);
assign cell_60_0 =
   (bitdata[227:227] == 1'b1 ? sw_0_0_13_down0 :
    bitdata[227:227] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[841:841] == 1'b1 ? sw_0_1_13_down0 :
    bitdata[841:841] == 1'b0 ? 1'b0 : 1'bx);
assign cell_61_0 =
   (bitdata[116:112] == 5'b11110 ? sw_0_0_8_down0 :
    bitdata[116:112] == 5'b00001 ? sw_0_0_8_down1 :
    bitdata[116:112] == 5'b10001 ? sw_0_0_8_down2 :
    bitdata[116:112] == 5'b01001 ? sw_0_0_8_down3 :
    bitdata[116:112] == 5'b11001 ? sw_0_0_8_down4 :
    bitdata[116:112] == 5'b10000 ? cell_71_5 :
    bitdata[116:112] == 5'b01000 ? cell_71_6 :
    bitdata[116:112] == 5'b11000 ? cell_71_7 :
    bitdata[116:112] == 5'b00100 ? cell_71_8 :
    bitdata[116:112] == 5'b10100 ? cell_80_6 :
    bitdata[116:112] == 5'b01100 ? cell_80_7 :
    bitdata[116:112] == 5'b11100 ? cell_80_8 :
    bitdata[116:112] == 5'b00010 ? cell_80_9 :
    bitdata[116:112] == 5'b10010 ? cell_80_10 :
    bitdata[116:112] == 5'b01010 ? cell_80_11 :
    bitdata[116:112] == 5'b11010 ? cell_80_12 :
    bitdata[116:112] == 5'b00110 ? cell_80_13 :
    bitdata[116:112] == 5'b10110 ? cell_80_14 :
    bitdata[116:112] == 5'b01110 ? cell_80_15 :
    bitdata[116:112] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[789:786] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[789:786] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[789:786] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[789:786] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[789:786] == 4'b1000 ? cell_63_8 :
    bitdata[789:786] == 4'b0100 ? cell_63_9 :
    bitdata[789:786] == 4'b1100 ? cell_71_5 :
    bitdata[789:786] == 4'b0010 ? cell_71_6 :
    bitdata[789:786] == 4'b1010 ? cell_71_7 :
    bitdata[789:786] == 4'b0110 ? cell_71_8 :
    bitdata[789:786] == 4'b1110 ? cell_83_0 :
    bitdata[789:786] == 4'b0 ? 1'b0 : 1'bx);
assign cell_61_1 =
   (bitdata[121:117] == 5'b11110 ? sw_0_0_8_down0 :
    bitdata[121:117] == 5'b00001 ? sw_0_0_8_down1 :
    bitdata[121:117] == 5'b10001 ? sw_0_0_8_down2 :
    bitdata[121:117] == 5'b01001 ? sw_0_0_8_down3 :
    bitdata[121:117] == 5'b11001 ? sw_0_0_8_down4 :
    bitdata[121:117] == 5'b10000 ? cell_71_5 :
    bitdata[121:117] == 5'b01000 ? cell_71_6 :
    bitdata[121:117] == 5'b11000 ? cell_71_7 :
    bitdata[121:117] == 5'b00100 ? cell_71_8 :
    bitdata[121:117] == 5'b10100 ? cell_80_6 :
    bitdata[121:117] == 5'b01100 ? cell_80_7 :
    bitdata[121:117] == 5'b11100 ? cell_80_8 :
    bitdata[121:117] == 5'b00010 ? cell_80_9 :
    bitdata[121:117] == 5'b10010 ? cell_80_10 :
    bitdata[121:117] == 5'b01010 ? cell_80_11 :
    bitdata[121:117] == 5'b11010 ? cell_80_12 :
    bitdata[121:117] == 5'b00110 ? cell_80_13 :
    bitdata[121:117] == 5'b10110 ? cell_80_14 :
    bitdata[121:117] == 5'b01110 ? cell_80_15 :
    bitdata[121:117] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[793:790] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[793:790] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[793:790] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[793:790] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[793:790] == 4'b1000 ? cell_63_8 :
    bitdata[793:790] == 4'b0100 ? cell_63_9 :
    bitdata[793:790] == 4'b1100 ? cell_71_5 :
    bitdata[793:790] == 4'b0010 ? cell_71_6 :
    bitdata[793:790] == 4'b1010 ? cell_71_7 :
    bitdata[793:790] == 4'b0110 ? cell_71_8 :
    bitdata[793:790] == 4'b1110 ? cell_83_0 :
    bitdata[793:790] == 4'b0 ? 1'b0 : 1'bx);
assign cell_61_2 =
   (bitdata[126:122] == 5'b11110 ? sw_0_0_8_down0 :
    bitdata[126:122] == 5'b00001 ? sw_0_0_8_down1 :
    bitdata[126:122] == 5'b10001 ? sw_0_0_8_down2 :
    bitdata[126:122] == 5'b01001 ? sw_0_0_8_down3 :
    bitdata[126:122] == 5'b11001 ? sw_0_0_8_down4 :
    bitdata[126:122] == 5'b10000 ? cell_71_5 :
    bitdata[126:122] == 5'b01000 ? cell_71_6 :
    bitdata[126:122] == 5'b11000 ? cell_71_7 :
    bitdata[126:122] == 5'b00100 ? cell_71_8 :
    bitdata[126:122] == 5'b10100 ? cell_80_6 :
    bitdata[126:122] == 5'b01100 ? cell_80_7 :
    bitdata[126:122] == 5'b11100 ? cell_80_8 :
    bitdata[126:122] == 5'b00010 ? cell_80_9 :
    bitdata[126:122] == 5'b10010 ? cell_80_10 :
    bitdata[126:122] == 5'b01010 ? cell_80_11 :
    bitdata[126:122] == 5'b11010 ? cell_80_12 :
    bitdata[126:122] == 5'b00110 ? cell_80_13 :
    bitdata[126:122] == 5'b10110 ? cell_80_14 :
    bitdata[126:122] == 5'b01110 ? cell_80_15 :
    bitdata[126:122] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[797:794] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[797:794] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[797:794] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[797:794] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[797:794] == 4'b1000 ? cell_63_8 :
    bitdata[797:794] == 4'b0100 ? cell_63_9 :
    bitdata[797:794] == 4'b1100 ? cell_71_5 :
    bitdata[797:794] == 4'b0010 ? cell_71_6 :
    bitdata[797:794] == 4'b1010 ? cell_71_7 :
    bitdata[797:794] == 4'b0110 ? cell_71_8 :
    bitdata[797:794] == 4'b1110 ? cell_83_0 :
    bitdata[797:794] == 4'b0 ? 1'b0 : 1'bx);
assign cell_61_3 =
   (bitdata[131:127] == 5'b11110 ? sw_0_0_8_down0 :
    bitdata[131:127] == 5'b00001 ? sw_0_0_8_down1 :
    bitdata[131:127] == 5'b10001 ? sw_0_0_8_down2 :
    bitdata[131:127] == 5'b01001 ? sw_0_0_8_down3 :
    bitdata[131:127] == 5'b11001 ? sw_0_0_8_down4 :
    bitdata[131:127] == 5'b10000 ? cell_71_5 :
    bitdata[131:127] == 5'b01000 ? cell_71_6 :
    bitdata[131:127] == 5'b11000 ? cell_71_7 :
    bitdata[131:127] == 5'b00100 ? cell_71_8 :
    bitdata[131:127] == 5'b10100 ? cell_80_6 :
    bitdata[131:127] == 5'b01100 ? cell_80_7 :
    bitdata[131:127] == 5'b11100 ? cell_80_8 :
    bitdata[131:127] == 5'b00010 ? cell_80_9 :
    bitdata[131:127] == 5'b10010 ? cell_80_10 :
    bitdata[131:127] == 5'b01010 ? cell_80_11 :
    bitdata[131:127] == 5'b11010 ? cell_80_12 :
    bitdata[131:127] == 5'b00110 ? cell_80_13 :
    bitdata[131:127] == 5'b10110 ? cell_80_14 :
    bitdata[131:127] == 5'b01110 ? cell_80_15 :
    bitdata[131:127] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[801:798] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[801:798] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[801:798] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[801:798] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[801:798] == 4'b1000 ? cell_63_8 :
    bitdata[801:798] == 4'b0100 ? cell_63_9 :
    bitdata[801:798] == 4'b1100 ? cell_71_5 :
    bitdata[801:798] == 4'b0010 ? cell_71_6 :
    bitdata[801:798] == 4'b1010 ? cell_71_7 :
    bitdata[801:798] == 4'b0110 ? cell_71_8 :
    bitdata[801:798] == 4'b1110 ? cell_83_0 :
    bitdata[801:798] == 4'b0 ? 1'b0 : 1'bx);
assign cell_61_4 =
   (bitdata[1064:1063] == 2'b11 ? sw_2_0_4_down0 :
    bitdata[1064:1063] == 2'b10 ? cell_79_3 :
    bitdata[1064:1063] == 2'b01 ? cell_91_0 :
    bitdata[1064:1063] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1200:1198] == 3'b001 ? sw_2_1_8_down0 :
    bitdata[1200:1198] == 3'b100 ? cell_62_5 :
    bitdata[1200:1198] == 3'b010 ? cell_64_6 :
    bitdata[1200:1198] == 3'b110 ? cell_64_7 :
    bitdata[1200:1198] == 3'b0 ? 16'b0 : 16'bx);
assign cell_62_0 =
   (bitdata[183:181] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[183:181] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[183:181] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[183:181] == 3'b100 ? cell_64_8 :
    bitdata[183:181] == 3'b010 ? cell_64_9 :
    bitdata[183:181] == 3'b110 ? cell_83_0 :
    bitdata[183:181] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[737:734] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[737:734] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[737:734] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[737:734] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[737:734] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[737:734] == 4'b1000 ? cell_64_8 :
    bitdata[737:734] == 4'b0100 ? cell_64_9 :
    bitdata[737:734] == 4'b1100 ? cell_82_0 :
    bitdata[737:734] == 4'b0 ? 1'b0 : 1'bx);
assign cell_62_1 =
   (bitdata[186:184] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[186:184] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[186:184] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[186:184] == 3'b100 ? cell_64_8 :
    bitdata[186:184] == 3'b010 ? cell_64_9 :
    bitdata[186:184] == 3'b110 ? cell_83_0 :
    bitdata[186:184] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[741:738] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[741:738] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[741:738] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[741:738] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[741:738] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[741:738] == 4'b1000 ? cell_64_8 :
    bitdata[741:738] == 4'b0100 ? cell_64_9 :
    bitdata[741:738] == 4'b1100 ? cell_82_0 :
    bitdata[741:738] == 4'b0 ? 1'b0 : 1'bx);
assign cell_62_2 =
   (bitdata[189:187] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[189:187] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[189:187] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[189:187] == 3'b100 ? cell_64_8 :
    bitdata[189:187] == 3'b010 ? cell_64_9 :
    bitdata[189:187] == 3'b110 ? cell_83_0 :
    bitdata[189:187] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[745:742] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[745:742] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[745:742] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[745:742] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[745:742] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[745:742] == 4'b1000 ? cell_64_8 :
    bitdata[745:742] == 4'b0100 ? cell_64_9 :
    bitdata[745:742] == 4'b1100 ? cell_82_0 :
    bitdata[745:742] == 4'b0 ? 1'b0 : 1'bx);
assign cell_62_3 =
   (bitdata[192:190] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[192:190] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[192:190] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[192:190] == 3'b100 ? cell_64_8 :
    bitdata[192:190] == 3'b010 ? cell_64_9 :
    bitdata[192:190] == 3'b110 ? cell_83_0 :
    bitdata[192:190] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[749:746] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[749:746] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[749:746] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[749:746] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[749:746] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[749:746] == 4'b1000 ? cell_64_8 :
    bitdata[749:746] == 4'b0100 ? cell_64_9 :
    bitdata[749:746] == 4'b1100 ? cell_82_0 :
    bitdata[749:746] == 4'b0 ? 1'b0 : 1'bx);
assign cell_62_4 =
   (bitdata[1054:1052] == 3'b101 ? sw_2_0_3_down0 :
    bitdata[1054:1052] == 3'b100 ? cell_63_6 :
    bitdata[1054:1052] == 3'b010 ? cell_63_7 :
    bitdata[1054:1052] == 3'b110 ? cell_93_0 :
    bitdata[1054:1052] == 3'b001 ? cell_94_0 :
    bitdata[1054:1052] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1203:1201] == 3'b001 ? sw_2_1_8_down0 :
    bitdata[1203:1201] == 3'b100 ? cell_61_5 :
    bitdata[1203:1201] == 3'b010 ? cell_64_6 :
    bitdata[1203:1201] == 3'b110 ? cell_64_7 :
    bitdata[1203:1201] == 3'b0 ? 16'b0 : 16'bx);
assign cell_63_0 =
   (bitdata[307:303] == 5'b00001 ? sw_0_0_25_down0 :
    bitdata[307:303] == 5'b10001 ? sw_0_0_25_down1 :
    bitdata[307:303] == 5'b01001 ? sw_0_0_25_down2 :
    bitdata[307:303] == 5'b10000 ? cell_81_10 :
    bitdata[307:303] == 5'b01000 ? cell_81_11 :
    bitdata[307:303] == 5'b11000 ? cell_81_12 :
    bitdata[307:303] == 5'b00100 ? cell_81_13 :
    bitdata[307:303] == 5'b10100 ? cell_81_14 :
    bitdata[307:303] == 5'b01100 ? cell_81_15 :
    bitdata[307:303] == 5'b11100 ? cell_81_16 :
    bitdata[307:303] == 5'b00010 ? cell_81_17 :
    bitdata[307:303] == 5'b10010 ? cell_81_18 :
    bitdata[307:303] == 5'b01010 ? cell_81_19 :
    bitdata[307:303] == 5'b11010 ? cell_81_20 :
    bitdata[307:303] == 5'b00110 ? cell_81_21 :
    bitdata[307:303] == 5'b10110 ? cell_81_22 :
    bitdata[307:303] == 5'b01110 ? cell_81_23 :
    bitdata[307:303] == 5'b11110 ? cell_81_24 :
    bitdata[307:303] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[805:802] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[805:802] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[805:802] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[805:802] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[805:802] == 4'b1000 ? cell_61_6 :
    bitdata[805:802] == 4'b0100 ? cell_61_7 :
    bitdata[805:802] == 4'b1100 ? cell_71_5 :
    bitdata[805:802] == 4'b0010 ? cell_71_6 :
    bitdata[805:802] == 4'b1010 ? cell_71_7 :
    bitdata[805:802] == 4'b0110 ? cell_71_8 :
    bitdata[805:802] == 4'b1110 ? cell_83_0 :
    bitdata[805:802] == 4'b0 ? 1'b0 : 1'bx);
assign cell_63_1 =
   (bitdata[312:308] == 5'b00001 ? sw_0_0_25_down0 :
    bitdata[312:308] == 5'b10001 ? sw_0_0_25_down1 :
    bitdata[312:308] == 5'b01001 ? sw_0_0_25_down2 :
    bitdata[312:308] == 5'b10000 ? cell_81_10 :
    bitdata[312:308] == 5'b01000 ? cell_81_11 :
    bitdata[312:308] == 5'b11000 ? cell_81_12 :
    bitdata[312:308] == 5'b00100 ? cell_81_13 :
    bitdata[312:308] == 5'b10100 ? cell_81_14 :
    bitdata[312:308] == 5'b01100 ? cell_81_15 :
    bitdata[312:308] == 5'b11100 ? cell_81_16 :
    bitdata[312:308] == 5'b00010 ? cell_81_17 :
    bitdata[312:308] == 5'b10010 ? cell_81_18 :
    bitdata[312:308] == 5'b01010 ? cell_81_19 :
    bitdata[312:308] == 5'b11010 ? cell_81_20 :
    bitdata[312:308] == 5'b00110 ? cell_81_21 :
    bitdata[312:308] == 5'b10110 ? cell_81_22 :
    bitdata[312:308] == 5'b01110 ? cell_81_23 :
    bitdata[312:308] == 5'b11110 ? cell_81_24 :
    bitdata[312:308] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[809:806] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[809:806] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[809:806] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[809:806] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[809:806] == 4'b1000 ? cell_61_6 :
    bitdata[809:806] == 4'b0100 ? cell_61_7 :
    bitdata[809:806] == 4'b1100 ? cell_71_5 :
    bitdata[809:806] == 4'b0010 ? cell_71_6 :
    bitdata[809:806] == 4'b1010 ? cell_71_7 :
    bitdata[809:806] == 4'b0110 ? cell_71_8 :
    bitdata[809:806] == 4'b1110 ? cell_83_0 :
    bitdata[809:806] == 4'b0 ? 1'b0 : 1'bx);
assign cell_63_2 =
   (bitdata[317:313] == 5'b00001 ? sw_0_0_25_down0 :
    bitdata[317:313] == 5'b10001 ? sw_0_0_25_down1 :
    bitdata[317:313] == 5'b01001 ? sw_0_0_25_down2 :
    bitdata[317:313] == 5'b10000 ? cell_81_10 :
    bitdata[317:313] == 5'b01000 ? cell_81_11 :
    bitdata[317:313] == 5'b11000 ? cell_81_12 :
    bitdata[317:313] == 5'b00100 ? cell_81_13 :
    bitdata[317:313] == 5'b10100 ? cell_81_14 :
    bitdata[317:313] == 5'b01100 ? cell_81_15 :
    bitdata[317:313] == 5'b11100 ? cell_81_16 :
    bitdata[317:313] == 5'b00010 ? cell_81_17 :
    bitdata[317:313] == 5'b10010 ? cell_81_18 :
    bitdata[317:313] == 5'b01010 ? cell_81_19 :
    bitdata[317:313] == 5'b11010 ? cell_81_20 :
    bitdata[317:313] == 5'b00110 ? cell_81_21 :
    bitdata[317:313] == 5'b10110 ? cell_81_22 :
    bitdata[317:313] == 5'b01110 ? cell_81_23 :
    bitdata[317:313] == 5'b11110 ? cell_81_24 :
    bitdata[317:313] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[813:810] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[813:810] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[813:810] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[813:810] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[813:810] == 4'b1000 ? cell_61_6 :
    bitdata[813:810] == 4'b0100 ? cell_61_7 :
    bitdata[813:810] == 4'b1100 ? cell_71_5 :
    bitdata[813:810] == 4'b0010 ? cell_71_6 :
    bitdata[813:810] == 4'b1010 ? cell_71_7 :
    bitdata[813:810] == 4'b0110 ? cell_71_8 :
    bitdata[813:810] == 4'b1110 ? cell_83_0 :
    bitdata[813:810] == 4'b0 ? 1'b0 : 1'bx);
assign cell_63_3 =
   (bitdata[322:318] == 5'b00001 ? sw_0_0_25_down0 :
    bitdata[322:318] == 5'b10001 ? sw_0_0_25_down1 :
    bitdata[322:318] == 5'b01001 ? sw_0_0_25_down2 :
    bitdata[322:318] == 5'b10000 ? cell_81_10 :
    bitdata[322:318] == 5'b01000 ? cell_81_11 :
    bitdata[322:318] == 5'b11000 ? cell_81_12 :
    bitdata[322:318] == 5'b00100 ? cell_81_13 :
    bitdata[322:318] == 5'b10100 ? cell_81_14 :
    bitdata[322:318] == 5'b01100 ? cell_81_15 :
    bitdata[322:318] == 5'b11100 ? cell_81_16 :
    bitdata[322:318] == 5'b00010 ? cell_81_17 :
    bitdata[322:318] == 5'b10010 ? cell_81_18 :
    bitdata[322:318] == 5'b01010 ? cell_81_19 :
    bitdata[322:318] == 5'b11010 ? cell_81_20 :
    bitdata[322:318] == 5'b00110 ? cell_81_21 :
    bitdata[322:318] == 5'b10110 ? cell_81_22 :
    bitdata[322:318] == 5'b01110 ? cell_81_23 :
    bitdata[322:318] == 5'b11110 ? cell_81_24 :
    bitdata[322:318] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[817:814] == 4'b0001 ? sw_0_1_11_down0 :
    bitdata[817:814] == 4'b1001 ? sw_0_1_11_down1 :
    bitdata[817:814] == 4'b0101 ? sw_0_1_11_down2 :
    bitdata[817:814] == 4'b1101 ? sw_0_1_11_down3 :
    bitdata[817:814] == 4'b1000 ? cell_61_6 :
    bitdata[817:814] == 4'b0100 ? cell_61_7 :
    bitdata[817:814] == 4'b1100 ? cell_71_5 :
    bitdata[817:814] == 4'b0010 ? cell_71_6 :
    bitdata[817:814] == 4'b1010 ? cell_71_7 :
    bitdata[817:814] == 4'b0110 ? cell_71_8 :
    bitdata[817:814] == 4'b1110 ? cell_83_0 :
    bitdata[817:814] == 4'b0 ? 1'b0 : 1'bx);
assign cell_63_4 =
   (bitdata[1057:1055] == 3'b001 ? sw_2_0_3_down0 :
    bitdata[1057:1055] == 3'b100 ? cell_62_5 :
    bitdata[1057:1055] == 3'b010 ? cell_93_0 :
    bitdata[1057:1055] == 3'b110 ? cell_94_0 :
    bitdata[1057:1055] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1159:1157] == 3'b001 ? sw_2_1_5_down0 :
    bitdata[1159:1157] == 3'b100 ? cell_79_3 :
    bitdata[1159:1157] == 3'b010 ? cell_90_0 :
    bitdata[1159:1157] == 3'b110 ? cell_91_0 :
    bitdata[1159:1157] == 3'b0 ? 16'b0 : 16'bx);
assign cell_63_5 =
   (bitdata[1060:1058] == 3'b001 ? sw_2_0_3_down0 :
    bitdata[1060:1058] == 3'b100 ? cell_62_5 :
    bitdata[1060:1058] == 3'b010 ? cell_93_0 :
    bitdata[1060:1058] == 3'b110 ? cell_94_0 :
    bitdata[1060:1058] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1162:1160] == 3'b001 ? sw_2_1_5_down0 :
    bitdata[1162:1160] == 3'b100 ? cell_79_3 :
    bitdata[1162:1160] == 3'b010 ? cell_90_0 :
    bitdata[1162:1160] == 3'b110 ? cell_91_0 :
    bitdata[1162:1160] == 3'b0 ? 16'b0 : 16'bx);
assign cell_64_0 =
   (bitdata[195:193] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[195:193] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[195:193] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[195:193] == 3'b100 ? cell_62_6 :
    bitdata[195:193] == 3'b010 ? cell_62_7 :
    bitdata[195:193] == 3'b110 ? cell_83_0 :
    bitdata[195:193] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[753:750] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[753:750] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[753:750] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[753:750] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[753:750] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[753:750] == 4'b1000 ? cell_62_6 :
    bitdata[753:750] == 4'b0100 ? cell_62_7 :
    bitdata[753:750] == 4'b1100 ? cell_82_0 :
    bitdata[753:750] == 4'b0 ? 1'b0 : 1'bx);
assign cell_64_1 =
   (bitdata[198:196] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[198:196] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[198:196] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[198:196] == 3'b100 ? cell_62_6 :
    bitdata[198:196] == 3'b010 ? cell_62_7 :
    bitdata[198:196] == 3'b110 ? cell_83_0 :
    bitdata[198:196] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[757:754] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[757:754] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[757:754] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[757:754] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[757:754] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[757:754] == 4'b1000 ? cell_62_6 :
    bitdata[757:754] == 4'b0100 ? cell_62_7 :
    bitdata[757:754] == 4'b1100 ? cell_82_0 :
    bitdata[757:754] == 4'b0 ? 1'b0 : 1'bx);
assign cell_64_2 =
   (bitdata[201:199] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[201:199] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[201:199] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[201:199] == 3'b100 ? cell_62_6 :
    bitdata[201:199] == 3'b010 ? cell_62_7 :
    bitdata[201:199] == 3'b110 ? cell_83_0 :
    bitdata[201:199] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[761:758] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[761:758] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[761:758] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[761:758] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[761:758] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[761:758] == 4'b1000 ? cell_62_6 :
    bitdata[761:758] == 4'b0100 ? cell_62_7 :
    bitdata[761:758] == 4'b1100 ? cell_82_0 :
    bitdata[761:758] == 4'b0 ? 1'b0 : 1'bx);
assign cell_64_3 =
   (bitdata[204:202] == 3'b001 ? sw_0_0_10_down0 :
    bitdata[204:202] == 3'b101 ? sw_0_0_10_down1 :
    bitdata[204:202] == 3'b011 ? sw_0_0_10_down2 :
    bitdata[204:202] == 3'b100 ? cell_62_6 :
    bitdata[204:202] == 3'b010 ? cell_62_7 :
    bitdata[204:202] == 3'b110 ? cell_83_0 :
    bitdata[204:202] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[765:762] == 4'b0010 ? sw_0_1_10_down0 :
    bitdata[765:762] == 4'b1010 ? sw_0_1_10_down1 :
    bitdata[765:762] == 4'b0110 ? sw_0_1_10_down2 :
    bitdata[765:762] == 4'b1110 ? sw_0_1_10_down3 :
    bitdata[765:762] == 4'b0001 ? sw_0_1_10_down4 :
    bitdata[765:762] == 4'b1000 ? cell_62_6 :
    bitdata[765:762] == 4'b0100 ? cell_62_7 :
    bitdata[765:762] == 4'b1100 ? cell_82_0 :
    bitdata[765:762] == 4'b0 ? 1'b0 : 1'bx);
assign cell_64_4 =
   (bitdata[1094:1092] == 3'b001 ? sw_2_0_6_down0 :
    bitdata[1094:1092] == 3'b100 ? cell_76_2 :
    bitdata[1094:1092] == 3'b010 ? cell_92_0 :
    bitdata[1094:1092] == 3'b110 ? cell_95_0 :
    bitdata[1094:1092] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1205:1204] == 2'b11 ? sw_2_1_8_down0 :
    bitdata[1205:1204] == 2'b10 ? cell_61_5 :
    bitdata[1205:1204] == 2'b01 ? cell_62_5 :
    bitdata[1205:1204] == 2'b0 ? 16'b0 : 16'bx);
assign cell_64_5 =
   (bitdata[1097:1095] == 3'b001 ? sw_2_0_6_down0 :
    bitdata[1097:1095] == 3'b100 ? cell_76_2 :
    bitdata[1097:1095] == 3'b010 ? cell_92_0 :
    bitdata[1097:1095] == 3'b110 ? cell_95_0 :
    bitdata[1097:1095] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1207:1206] == 2'b11 ? sw_2_1_8_down0 :
    bitdata[1207:1206] == 2'b10 ? cell_61_5 :
    bitdata[1207:1206] == 2'b01 ? cell_62_5 :
    bitdata[1207:1206] == 2'b0 ? 16'b0 : 16'bx);
assign cell_65_0 =
   (bitdata[1101:1100] == 2'b11 ? sw_2_0_7_down0 :
    bitdata[1101:1100] == 2'b10 ? cell_66_1 :
    bitdata[1101:1100] == 2'b01 ? cell_71_3 :
    bitdata[1101:1100] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1189:1187] == 3'b001 ? sw_2_1_7_down0 :
    bitdata[1189:1187] == 3'b101 ? sw_2_1_7_down1 :
    bitdata[1189:1187] == 3'b100 ? cell_2_0 :
    bitdata[1189:1187] == 3'b010 ? cell_66_1 :
    bitdata[1189:1187] == 3'b110 ? cell_76_2 :
    bitdata[1189:1187] == 3'b0 ? 16'b0 : 16'bx);
assign cell_65_1 =
   (bitdata[1103:1102] == 2'b11 ? sw_2_0_7_down0 :
    bitdata[1103:1102] == 2'b10 ? cell_66_1 :
    bitdata[1103:1102] == 2'b01 ? cell_71_3 :
    bitdata[1103:1102] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1192:1190] == 3'b001 ? sw_2_1_7_down0 :
    bitdata[1192:1190] == 3'b101 ? sw_2_1_7_down1 :
    bitdata[1192:1190] == 3'b100 ? cell_2_0 :
    bitdata[1192:1190] == 3'b010 ? cell_66_1 :
    bitdata[1192:1190] == 3'b110 ? cell_76_2 :
    bitdata[1192:1190] == 3'b0 ? 16'b0 : 16'bx);
assign cell_66_0 =
   (bitdata[1105:1104] == 2'b11 ? sw_2_0_7_down0 :
    bitdata[1105:1104] == 2'b10 ? cell_65_2 :
    bitdata[1105:1104] == 2'b01 ? cell_71_3 :
    bitdata[1105:1104] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1195:1193] == 3'b001 ? sw_2_1_7_down0 :
    bitdata[1195:1193] == 3'b101 ? sw_2_1_7_down1 :
    bitdata[1195:1193] == 3'b100 ? cell_2_0 :
    bitdata[1195:1193] == 3'b010 ? cell_65_2 :
    bitdata[1195:1193] == 3'b110 ? cell_76_2 :
    bitdata[1195:1193] == 3'b0 ? 16'b0 : 16'bx);
assign cell_66_2 =
   (bitdata[216:214] == 3'b011 ? sw_0_0_12_down0 :
    bitdata[216:214] == 3'b100 ? cell_8_0 :
    bitdata[216:214] == 3'b010 ? cell_72_5 :
    bitdata[216:214] == 3'b110 ? cell_72_6 :
    bitdata[216:214] == 3'b001 ? cell_72_7 :
    bitdata[216:214] == 3'b101 ? cell_72_8 :
    bitdata[216:214] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[630:626] == 5'b01011 ? sw_0_1_8_down0 :
    bitdata[630:626] == 5'b11011 ? sw_0_1_8_down1 :
    bitdata[630:626] == 5'b00111 ? sw_0_1_8_down2 :
    bitdata[630:626] == 5'b10111 ? sw_0_1_8_down3 :
    bitdata[630:626] == 5'b01111 ? sw_0_1_8_down4 :
    bitdata[630:626] == 5'b11111 ? sw_0_1_8_down5 :
    bitdata[630:626] == 5'b10000 ? cell_80_6 :
    bitdata[630:626] == 5'b01000 ? cell_80_7 :
    bitdata[630:626] == 5'b11000 ? cell_80_8 :
    bitdata[630:626] == 5'b00100 ? cell_80_9 :
    bitdata[630:626] == 5'b10100 ? cell_80_10 :
    bitdata[630:626] == 5'b01100 ? cell_80_11 :
    bitdata[630:626] == 5'b11100 ? cell_80_12 :
    bitdata[630:626] == 5'b00010 ? cell_80_13 :
    bitdata[630:626] == 5'b10010 ? cell_80_14 :
    bitdata[630:626] == 5'b01010 ? cell_80_15 :
    bitdata[630:626] == 5'b11010 ? cell_81_10 :
    bitdata[630:626] == 5'b00110 ? cell_81_11 :
    bitdata[630:626] == 5'b10110 ? cell_81_12 :
    bitdata[630:626] == 5'b01110 ? cell_81_13 :
    bitdata[630:626] == 5'b11110 ? cell_81_14 :
    bitdata[630:626] == 5'b00001 ? cell_81_15 :
    bitdata[630:626] == 5'b10001 ? cell_81_16 :
    bitdata[630:626] == 5'b01001 ? cell_81_17 :
    bitdata[630:626] == 5'b11001 ? cell_81_18 :
    bitdata[630:626] == 5'b00101 ? cell_81_19 :
    bitdata[630:626] == 5'b10101 ? cell_81_20 :
    bitdata[630:626] == 5'b01101 ? cell_81_21 :
    bitdata[630:626] == 5'b11101 ? cell_81_22 :
    bitdata[630:626] == 5'b00011 ? cell_81_23 :
    bitdata[630:626] == 5'b10011 ? cell_81_24 :
    bitdata[630:626] == 5'b0 ? 1'b0 : 1'bx);
assign cell_67_0 =
   (bitdata[1076:1074] == 3'b001 ? sw_2_0_5_down0 :
    bitdata[1076:1074] == 3'b100 ? cell_72_3 :
    bitdata[1076:1074] == 3'b010 ? cell_77_2 :
    bitdata[1076:1074] == 3'b110 ? cell_78_3 :
    bitdata[1076:1074] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1175:1173] == 3'b001 ? sw_2_1_6_down0 :
    bitdata[1175:1173] == 3'b100 ? cell_68_1 :
    bitdata[1175:1173] == 3'b010 ? cell_72_3 :
    bitdata[1175:1173] == 3'b110 ? cell_77_2 :
    bitdata[1175:1173] == 3'b0 ? 16'b0 : 16'bx);
assign cell_67_2 =
   (bitdata[240:240] == 1'b1 ? sw_0_0_17_down0 :
    bitdata[240:240] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[827:826] == 2'b10 ? sw_0_1_12_down0 :
    bitdata[827:826] == 2'b01 ? sw_0_1_12_down1 :
    bitdata[827:826] == 2'b0 ? 1'b0 : 1'bx);
assign cell_68_0 =
   (bitdata[1116:1115] == 2'b11 ? sw_2_0_8_down0 :
    bitdata[1116:1115] == 2'b10 ? cell_2_0 :
    bitdata[1116:1115] == 2'b01 ? cell_90_0 :
    bitdata[1116:1115] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1178:1176] == 3'b001 ? sw_2_1_6_down0 :
    bitdata[1178:1176] == 3'b100 ? cell_67_1 :
    bitdata[1178:1176] == 3'b010 ? cell_72_3 :
    bitdata[1178:1176] == 3'b110 ? cell_77_2 :
    bitdata[1178:1176] == 3'b0 ? 16'b0 : 16'bx);
assign cell_68_2 =
   (bitdata[241:241] == 1'b1 ? sw_0_0_17_down0 :
    bitdata[241:241] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[829:828] == 2'b10 ? sw_0_1_12_down0 :
    bitdata[829:828] == 2'b01 ? sw_0_1_12_down1 :
    bitdata[829:828] == 2'b0 ? 1'b0 : 1'bx);
assign cell_69_0 =
   (bitdata[960:959] == 2'b01 ? sw_1_0_6_down0 :
    bitdata[960:959] == 2'b10 ? cell_70_1 :
    bitdata[960:959] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[1026:1024] == 3'b001 ? sw_1_1_6_down0 :
    bitdata[1026:1024] == 3'b100 ? cell_5_0 :
    bitdata[1026:1024] == 3'b010 ? cell_38_0 :
    bitdata[1026:1024] == 3'b110 ? cell_70_1 :
    bitdata[1026:1024] == 3'b0 ? 8'b0 : 8'bx);
assign cell_69_2 =
   (bitdata[261:261] == 1'b1 ? sw_0_0_21_down0 :
    bitdata[261:261] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[635:631] == 5'b01011 ? sw_0_1_8_down0 :
    bitdata[635:631] == 5'b11011 ? sw_0_1_8_down1 :
    bitdata[635:631] == 5'b00111 ? sw_0_1_8_down2 :
    bitdata[635:631] == 5'b10111 ? sw_0_1_8_down3 :
    bitdata[635:631] == 5'b01111 ? sw_0_1_8_down4 :
    bitdata[635:631] == 5'b11111 ? sw_0_1_8_down5 :
    bitdata[635:631] == 5'b10000 ? cell_80_6 :
    bitdata[635:631] == 5'b01000 ? cell_80_7 :
    bitdata[635:631] == 5'b11000 ? cell_80_8 :
    bitdata[635:631] == 5'b00100 ? cell_80_9 :
    bitdata[635:631] == 5'b10100 ? cell_80_10 :
    bitdata[635:631] == 5'b01100 ? cell_80_11 :
    bitdata[635:631] == 5'b11100 ? cell_80_12 :
    bitdata[635:631] == 5'b00010 ? cell_80_13 :
    bitdata[635:631] == 5'b10010 ? cell_80_14 :
    bitdata[635:631] == 5'b01010 ? cell_80_15 :
    bitdata[635:631] == 5'b11010 ? cell_81_10 :
    bitdata[635:631] == 5'b00110 ? cell_81_11 :
    bitdata[635:631] == 5'b10110 ? cell_81_12 :
    bitdata[635:631] == 5'b01110 ? cell_81_13 :
    bitdata[635:631] == 5'b11110 ? cell_81_14 :
    bitdata[635:631] == 5'b00001 ? cell_81_15 :
    bitdata[635:631] == 5'b10001 ? cell_81_16 :
    bitdata[635:631] == 5'b01001 ? cell_81_17 :
    bitdata[635:631] == 5'b11001 ? cell_81_18 :
    bitdata[635:631] == 5'b00101 ? cell_81_19 :
    bitdata[635:631] == 5'b10101 ? cell_81_20 :
    bitdata[635:631] == 5'b01101 ? cell_81_21 :
    bitdata[635:631] == 5'b11101 ? cell_81_22 :
    bitdata[635:631] == 5'b00011 ? cell_81_23 :
    bitdata[635:631] == 5'b10011 ? cell_81_24 :
    bitdata[635:631] == 5'b0 ? 1'b0 : 1'bx);
assign cell_70_0 =
   (bitdata[962:961] == 2'b01 ? sw_1_0_6_down0 :
    bitdata[962:961] == 2'b10 ? cell_69_1 :
    bitdata[962:961] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[1029:1027] == 3'b001 ? sw_1_1_6_down0 :
    bitdata[1029:1027] == 3'b100 ? cell_5_0 :
    bitdata[1029:1027] == 3'b010 ? cell_38_0 :
    bitdata[1029:1027] == 3'b110 ? cell_69_1 :
    bitdata[1029:1027] == 3'b0 ? 8'b0 : 8'bx);
assign cell_70_2 =
   (bitdata[266:264] == 3'b001 ? sw_0_0_22_down0 :
    bitdata[266:264] == 3'b100 ? cell_19_0 :
    bitdata[266:264] == 3'b010 ? cell_20_0 :
    bitdata[266:264] == 3'b110 ? cell_21_0 :
    bitdata[266:264] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[769:766] == 4'b0110 ? sw_0_1_10_down0 :
    bitdata[769:766] == 4'b1110 ? sw_0_1_10_down1 :
    bitdata[769:766] == 4'b0001 ? sw_0_1_10_down2 :
    bitdata[769:766] == 4'b1001 ? sw_0_1_10_down3 :
    bitdata[769:766] == 4'b0101 ? sw_0_1_10_down4 :
    bitdata[769:766] == 4'b1000 ? cell_62_6 :
    bitdata[769:766] == 4'b0100 ? cell_62_7 :
    bitdata[769:766] == 4'b1100 ? cell_64_8 :
    bitdata[769:766] == 4'b0010 ? cell_64_9 :
    bitdata[769:766] == 4'b1010 ? cell_82_0 :
    bitdata[769:766] == 4'b0 ? 1'b0 : 1'bx);
assign cell_71_0 =
   (bitdata[136:132] == 5'b10110 ? sw_0_0_8_down0 :
    bitdata[136:132] == 5'b01110 ? sw_0_0_8_down1 :
    bitdata[136:132] == 5'b11110 ? sw_0_0_8_down2 :
    bitdata[136:132] == 5'b00001 ? sw_0_0_8_down3 :
    bitdata[136:132] == 5'b10001 ? sw_0_0_8_down4 :
    bitdata[136:132] == 5'b10000 ? cell_61_6 :
    bitdata[136:132] == 5'b01000 ? cell_61_7 :
    bitdata[136:132] == 5'b11000 ? cell_80_6 :
    bitdata[136:132] == 5'b00100 ? cell_80_7 :
    bitdata[136:132] == 5'b10100 ? cell_80_8 :
    bitdata[136:132] == 5'b01100 ? cell_80_9 :
    bitdata[136:132] == 5'b11100 ? cell_80_10 :
    bitdata[136:132] == 5'b00010 ? cell_80_11 :
    bitdata[136:132] == 5'b10010 ? cell_80_12 :
    bitdata[136:132] == 5'b01010 ? cell_80_13 :
    bitdata[136:132] == 5'b11010 ? cell_80_14 :
    bitdata[136:132] == 5'b00110 ? cell_80_15 :
    bitdata[136:132] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[821:818] == 4'b0110 ? sw_0_1_11_down0 :
    bitdata[821:818] == 4'b1110 ? sw_0_1_11_down1 :
    bitdata[821:818] == 4'b0001 ? sw_0_1_11_down2 :
    bitdata[821:818] == 4'b1001 ? sw_0_1_11_down3 :
    bitdata[821:818] == 4'b1000 ? cell_61_6 :
    bitdata[821:818] == 4'b0100 ? cell_61_7 :
    bitdata[821:818] == 4'b1100 ? cell_63_8 :
    bitdata[821:818] == 4'b0010 ? cell_63_9 :
    bitdata[821:818] == 4'b1010 ? cell_83_0 :
    bitdata[821:818] == 4'b0 ? 1'b0 : 1'bx);
assign cell_71_1 =
   (bitdata[1107:1106] == 2'b11 ? sw_2_0_7_down0 :
    bitdata[1107:1106] == 2'b10 ? cell_65_2 :
    bitdata[1107:1106] == 2'b01 ? cell_66_1 :
    bitdata[1107:1106] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1144:1142] == 3'b001 ? sw_2_1_4_down0 :
    bitdata[1144:1142] == 3'b100 ? cell_78_3 :
    bitdata[1144:1142] == 3'b010 ? cell_92_0 :
    bitdata[1144:1142] == 3'b110 ? cell_93_0 :
    bitdata[1144:1142] == 3'b0 ? 16'b0 : 16'bx);
assign cell_71_2 =
   (bitdata[1109:1108] == 2'b11 ? sw_2_0_7_down0 :
    bitdata[1109:1108] == 2'b10 ? cell_65_2 :
    bitdata[1109:1108] == 2'b01 ? cell_66_1 :
    bitdata[1109:1108] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1147:1145] == 3'b001 ? sw_2_1_4_down0 :
    bitdata[1147:1145] == 3'b100 ? cell_78_3 :
    bitdata[1147:1145] == 3'b010 ? cell_92_0 :
    bitdata[1147:1145] == 3'b110 ? cell_93_0 :
    bitdata[1147:1145] == 3'b0 ? 16'b0 : 16'bx);
assign cell_71_4 =
   (bitdata[141:137] == 5'b10110 ? sw_0_0_8_down0 :
    bitdata[141:137] == 5'b01110 ? sw_0_0_8_down1 :
    bitdata[141:137] == 5'b11110 ? sw_0_0_8_down2 :
    bitdata[141:137] == 5'b00001 ? sw_0_0_8_down3 :
    bitdata[141:137] == 5'b10001 ? sw_0_0_8_down4 :
    bitdata[141:137] == 5'b10000 ? cell_61_6 :
    bitdata[141:137] == 5'b01000 ? cell_61_7 :
    bitdata[141:137] == 5'b11000 ? cell_80_6 :
    bitdata[141:137] == 5'b00100 ? cell_80_7 :
    bitdata[141:137] == 5'b10100 ? cell_80_8 :
    bitdata[141:137] == 5'b01100 ? cell_80_9 :
    bitdata[141:137] == 5'b11100 ? cell_80_10 :
    bitdata[141:137] == 5'b00010 ? cell_80_11 :
    bitdata[141:137] == 5'b10010 ? cell_80_12 :
    bitdata[141:137] == 5'b01010 ? cell_80_13 :
    bitdata[141:137] == 5'b11010 ? cell_80_14 :
    bitdata[141:137] == 5'b00110 ? cell_80_15 :
    bitdata[141:137] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[825:822] == 4'b0110 ? sw_0_1_11_down0 :
    bitdata[825:822] == 4'b1110 ? sw_0_1_11_down1 :
    bitdata[825:822] == 4'b0001 ? sw_0_1_11_down2 :
    bitdata[825:822] == 4'b1001 ? sw_0_1_11_down3 :
    bitdata[825:822] == 4'b1000 ? cell_61_6 :
    bitdata[825:822] == 4'b0100 ? cell_61_7 :
    bitdata[825:822] == 4'b1100 ? cell_63_8 :
    bitdata[825:822] == 4'b0010 ? cell_63_9 :
    bitdata[825:822] == 4'b1010 ? cell_83_0 :
    bitdata[825:822] == 4'b0 ? 1'b0 : 1'bx);
assign cell_72_0 =
   (bitdata[218:217] == 2'b01 ? sw_0_0_12_down0 :
    bitdata[218:217] == 2'b10 ? cell_8_0 :
    bitdata[218:217] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[873:872] == 2'b10 ? sw_0_1_18_down0 :
    bitdata[873:872] == 2'b01 ? sw_0_1_18_down1 :
    bitdata[873:872] == 2'b11 ? sw_0_1_18_down2 :
    bitdata[873:872] == 2'b0 ? 1'b0 : 1'bx);
assign cell_72_1 =
   (bitdata[1079:1077] == 3'b001 ? sw_2_0_5_down0 :
    bitdata[1079:1077] == 3'b100 ? cell_67_1 :
    bitdata[1079:1077] == 3'b010 ? cell_77_2 :
    bitdata[1079:1077] == 3'b110 ? cell_78_3 :
    bitdata[1079:1077] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1181:1179] == 3'b001 ? sw_2_1_6_down0 :
    bitdata[1181:1179] == 3'b100 ? cell_67_1 :
    bitdata[1181:1179] == 3'b010 ? cell_68_1 :
    bitdata[1181:1179] == 3'b110 ? cell_77_2 :
    bitdata[1181:1179] == 3'b0 ? 16'b0 : 16'bx);
assign cell_72_2 =
   (bitdata[1082:1080] == 3'b001 ? sw_2_0_5_down0 :
    bitdata[1082:1080] == 3'b100 ? cell_67_1 :
    bitdata[1082:1080] == 3'b010 ? cell_77_2 :
    bitdata[1082:1080] == 3'b110 ? cell_78_3 :
    bitdata[1082:1080] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1184:1182] == 3'b001 ? sw_2_1_6_down0 :
    bitdata[1184:1182] == 3'b100 ? cell_67_1 :
    bitdata[1184:1182] == 3'b010 ? cell_68_1 :
    bitdata[1184:1182] == 3'b110 ? cell_77_2 :
    bitdata[1184:1182] == 3'b0 ? 16'b0 : 16'bx);
assign cell_72_4 =
   (bitdata[220:219] == 2'b01 ? sw_0_0_12_down0 :
    bitdata[220:219] == 2'b10 ? cell_8_0 :
    bitdata[220:219] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[875:874] == 2'b10 ? sw_0_1_18_down0 :
    bitdata[875:874] == 2'b01 ? sw_0_1_18_down1 :
    bitdata[875:874] == 2'b11 ? sw_0_1_18_down2 :
    bitdata[875:874] == 2'b0 ? 1'b0 : 1'bx);
assign cell_73_0 =
   (bitdata[930:928] == 3'b110 ? sw_1_0_3_down0 :
    bitdata[930:928] == 3'b001 ? sw_1_0_3_down1 :
    bitdata[930:928] == 3'b100 ? cell_87_0 :
    bitdata[930:928] == 3'b010 ? cell_89_0 :
    bitdata[930:928] == 3'b0 ? 8'b0 : 8'bx) |
   (bitdata[1006:1004] == 3'b110 ? sw_1_1_5_down0 :
    bitdata[1006:1004] == 3'b001 ? sw_1_1_5_down1 :
    bitdata[1006:1004] == 3'b100 ? cell_75_3 :
    bitdata[1006:1004] == 3'b010 ? cell_88_0 :
    bitdata[1006:1004] == 3'b0 ? 8'b0 : 8'bx);
assign cell_73_1 =
   (bitdata[933:931] == 3'b110 ? sw_1_0_3_down0 :
    bitdata[933:931] == 3'b001 ? sw_1_0_3_down1 :
    bitdata[933:931] == 3'b100 ? cell_87_0 :
    bitdata[933:931] == 3'b010 ? cell_89_0 :
    bitdata[933:931] == 3'b0 ? 8'b0 : 8'bx) |
   (bitdata[1009:1007] == 3'b110 ? sw_1_1_5_down0 :
    bitdata[1009:1007] == 3'b001 ? sw_1_1_5_down1 :
    bitdata[1009:1007] == 3'b100 ? cell_75_3 :
    bitdata[1009:1007] == 3'b010 ? cell_88_0 :
    bitdata[1009:1007] == 3'b0 ? 8'b0 : 8'bx);
assign cell_73_2 =
   (bitdata[936:934] == 3'b110 ? sw_1_0_3_down0 :
    bitdata[936:934] == 3'b001 ? sw_1_0_3_down1 :
    bitdata[936:934] == 3'b100 ? cell_87_0 :
    bitdata[936:934] == 3'b010 ? cell_89_0 :
    bitdata[936:934] == 3'b0 ? 8'b0 : 8'bx) |
   (bitdata[1012:1010] == 3'b110 ? sw_1_1_5_down0 :
    bitdata[1012:1010] == 3'b001 ? sw_1_1_5_down1 :
    bitdata[1012:1010] == 3'b100 ? cell_75_3 :
    bitdata[1012:1010] == 3'b010 ? cell_88_0 :
    bitdata[1012:1010] == 3'b0 ? 8'b0 : 8'bx);
assign cell_73_3 =
   (bitdata[939:937] == 3'b110 ? sw_1_0_3_down0 :
    bitdata[939:937] == 3'b001 ? sw_1_0_3_down1 :
    bitdata[939:937] == 3'b100 ? cell_87_0 :
    bitdata[939:937] == 3'b010 ? cell_89_0 :
    bitdata[939:937] == 3'b0 ? 8'b0 : 8'bx) |
   (bitdata[1015:1013] == 3'b110 ? sw_1_1_5_down0 :
    bitdata[1015:1013] == 3'b001 ? sw_1_1_5_down1 :
    bitdata[1015:1013] == 3'b100 ? cell_75_3 :
    bitdata[1015:1013] == 3'b010 ? cell_88_0 :
    bitdata[1015:1013] == 3'b0 ? 8'b0 : 8'bx);
assign cell_73_4 =
   (bitdata[327:323] == 5'b01001 ? sw_0_0_25_down0 :
    bitdata[327:323] == 5'b11001 ? sw_0_0_25_down1 :
    bitdata[327:323] == 5'b00101 ? sw_0_0_25_down2 :
    bitdata[327:323] == 5'b10000 ? cell_63_8 :
    bitdata[327:323] == 5'b01000 ? cell_63_9 :
    bitdata[327:323] == 5'b11000 ? cell_81_10 :
    bitdata[327:323] == 5'b00100 ? cell_81_11 :
    bitdata[327:323] == 5'b10100 ? cell_81_12 :
    bitdata[327:323] == 5'b01100 ? cell_81_13 :
    bitdata[327:323] == 5'b11100 ? cell_81_14 :
    bitdata[327:323] == 5'b00010 ? cell_81_15 :
    bitdata[327:323] == 5'b10010 ? cell_81_16 :
    bitdata[327:323] == 5'b01010 ? cell_81_17 :
    bitdata[327:323] == 5'b11010 ? cell_81_18 :
    bitdata[327:323] == 5'b00110 ? cell_81_19 :
    bitdata[327:323] == 5'b10110 ? cell_81_20 :
    bitdata[327:323] == 5'b01110 ? cell_81_21 :
    bitdata[327:323] == 5'b11110 ? cell_81_22 :
    bitdata[327:323] == 5'b00001 ? cell_81_23 :
    bitdata[327:323] == 5'b10001 ? cell_81_24 :
    bitdata[327:323] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[831:830] == 2'b10 ? sw_0_1_12_down0 :
    bitdata[831:830] == 2'b01 ? sw_0_1_12_down1 :
    bitdata[831:830] == 2'b0 ? 1'b0 : 1'bx);
assign cell_73_5 =
   (bitdata[332:328] == 5'b01001 ? sw_0_0_25_down0 :
    bitdata[332:328] == 5'b11001 ? sw_0_0_25_down1 :
    bitdata[332:328] == 5'b00101 ? sw_0_0_25_down2 :
    bitdata[332:328] == 5'b10000 ? cell_63_8 :
    bitdata[332:328] == 5'b01000 ? cell_63_9 :
    bitdata[332:328] == 5'b11000 ? cell_81_10 :
    bitdata[332:328] == 5'b00100 ? cell_81_11 :
    bitdata[332:328] == 5'b10100 ? cell_81_12 :
    bitdata[332:328] == 5'b01100 ? cell_81_13 :
    bitdata[332:328] == 5'b11100 ? cell_81_14 :
    bitdata[332:328] == 5'b00010 ? cell_81_15 :
    bitdata[332:328] == 5'b10010 ? cell_81_16 :
    bitdata[332:328] == 5'b01010 ? cell_81_17 :
    bitdata[332:328] == 5'b11010 ? cell_81_18 :
    bitdata[332:328] == 5'b00110 ? cell_81_19 :
    bitdata[332:328] == 5'b10110 ? cell_81_20 :
    bitdata[332:328] == 5'b01110 ? cell_81_21 :
    bitdata[332:328] == 5'b11110 ? cell_81_22 :
    bitdata[332:328] == 5'b00001 ? cell_81_23 :
    bitdata[332:328] == 5'b10001 ? cell_81_24 :
    bitdata[332:328] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[833:832] == 2'b10 ? sw_0_1_12_down0 :
    bitdata[833:832] == 2'b01 ? sw_0_1_12_down1 :
    bitdata[833:832] == 2'b0 ? 1'b0 : 1'bx);
assign cell_73_6 =
   (bitdata[337:333] == 5'b01001 ? sw_0_0_25_down0 :
    bitdata[337:333] == 5'b11001 ? sw_0_0_25_down1 :
    bitdata[337:333] == 5'b00101 ? sw_0_0_25_down2 :
    bitdata[337:333] == 5'b10000 ? cell_63_8 :
    bitdata[337:333] == 5'b01000 ? cell_63_9 :
    bitdata[337:333] == 5'b11000 ? cell_81_10 :
    bitdata[337:333] == 5'b00100 ? cell_81_11 :
    bitdata[337:333] == 5'b10100 ? cell_81_12 :
    bitdata[337:333] == 5'b01100 ? cell_81_13 :
    bitdata[337:333] == 5'b11100 ? cell_81_14 :
    bitdata[337:333] == 5'b00010 ? cell_81_15 :
    bitdata[337:333] == 5'b10010 ? cell_81_16 :
    bitdata[337:333] == 5'b01010 ? cell_81_17 :
    bitdata[337:333] == 5'b11010 ? cell_81_18 :
    bitdata[337:333] == 5'b00110 ? cell_81_19 :
    bitdata[337:333] == 5'b10110 ? cell_81_20 :
    bitdata[337:333] == 5'b01110 ? cell_81_21 :
    bitdata[337:333] == 5'b11110 ? cell_81_22 :
    bitdata[337:333] == 5'b00001 ? cell_81_23 :
    bitdata[337:333] == 5'b10001 ? cell_81_24 :
    bitdata[337:333] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[835:834] == 2'b10 ? sw_0_1_12_down0 :
    bitdata[835:834] == 2'b01 ? sw_0_1_12_down1 :
    bitdata[835:834] == 2'b0 ? 1'b0 : 1'bx);
assign cell_74_0 =
   (bitdata[948:947] == 2'b11 ? sw_1_0_4_down0 :
    bitdata[948:947] == 2'b10 ? cell_84_0 :
    bitdata[948:947] == 2'b01 ? cell_85_0 :
    bitdata[948:947] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[988:986] == 3'b001 ? sw_1_1_3_down0 :
    bitdata[988:986] == 3'b100 ? cell_86_0 :
    bitdata[988:986] == 3'b010 ? cell_87_0 :
    bitdata[988:986] == 3'b110 ? cell_89_0 :
    bitdata[988:986] == 3'b0 ? 8'b0 : 8'bx);
assign cell_74_1 =
   (bitdata[950:949] == 2'b11 ? sw_1_0_4_down0 :
    bitdata[950:949] == 2'b10 ? cell_84_0 :
    bitdata[950:949] == 2'b01 ? cell_85_0 :
    bitdata[950:949] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[991:989] == 3'b001 ? sw_1_1_3_down0 :
    bitdata[991:989] == 3'b100 ? cell_86_0 :
    bitdata[991:989] == 3'b010 ? cell_87_0 :
    bitdata[991:989] == 3'b110 ? cell_89_0 :
    bitdata[991:989] == 3'b0 ? 8'b0 : 8'bx);
assign cell_74_2 =
   (bitdata[371:370] == 2'b01 ? sw_0_0_26_down0 :
    bitdata[371:370] == 2'b11 ? sw_0_0_26_down1 :
    bitdata[371:370] == 2'b10 ? cell_6_0 :
    bitdata[371:370] == 2'b0 ? 1'b0 : 1'bx) |
   (bitdata[837:836] == 2'b10 ? sw_0_1_12_down0 :
    bitdata[837:836] == 2'b01 ? sw_0_1_12_down1 :
    bitdata[837:836] == 2'b0 ? 1'b0 : 1'bx);
assign cell_75_0 =
   (bitdata[955:954] == 2'b01 ? sw_1_0_5_down0 :
    bitdata[955:954] == 2'b10 ? cell_86_0 :
    bitdata[955:954] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[1018:1016] == 3'b110 ? sw_1_1_5_down0 :
    bitdata[1018:1016] == 3'b001 ? sw_1_1_5_down1 :
    bitdata[1018:1016] == 3'b100 ? cell_73_7 :
    bitdata[1018:1016] == 3'b010 ? cell_88_0 :
    bitdata[1018:1016] == 3'b0 ? 8'b0 : 8'bx);
assign cell_75_1 =
   (bitdata[957:956] == 2'b01 ? sw_1_0_5_down0 :
    bitdata[957:956] == 2'b10 ? cell_86_0 :
    bitdata[957:956] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[1021:1019] == 3'b110 ? sw_1_1_5_down0 :
    bitdata[1021:1019] == 3'b001 ? sw_1_1_5_down1 :
    bitdata[1021:1019] == 3'b100 ? cell_73_7 :
    bitdata[1021:1019] == 3'b010 ? cell_88_0 :
    bitdata[1021:1019] == 3'b0 ? 8'b0 : 8'bx);
assign cell_75_2 =
   (bitdata[223:221] == 3'b011 ? sw_0_0_12_down0 :
    bitdata[223:221] == 3'b100 ? cell_8_0 :
    bitdata[223:221] == 3'b010 ? cell_72_5 :
    bitdata[223:221] == 3'b110 ? cell_72_6 :
    bitdata[223:221] == 3'b001 ? cell_72_7 :
    bitdata[223:221] == 3'b101 ? cell_72_8 :
    bitdata[223:221] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[724:722] == 3'b010 ? sw_0_1_9_down0 :
    bitdata[724:722] == 3'b110 ? sw_0_1_9_down1 :
    bitdata[724:722] == 3'b001 ? sw_0_1_9_down2 :
    bitdata[724:722] == 3'b100 ? cell_43_0 :
    bitdata[724:722] == 3'b0 ? 1'b0 : 1'bx);
assign cell_76_0 =
   (bitdata[964:963] == 2'b11 ? sw_1_0_6_down0 :
    bitdata[964:963] == 2'b10 ? cell_69_1 :
    bitdata[964:963] == 2'b01 ? cell_70_1 :
    bitdata[964:963] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[995:994] == 2'b11 ? sw_1_1_4_down0 :
    bitdata[995:994] == 2'b10 ? cell_84_0 :
    bitdata[995:994] == 2'b01 ? cell_85_0 :
    bitdata[995:994] == 2'b0 ? 8'b0 : 8'bx);
assign cell_76_1 =
   (bitdata[966:965] == 2'b11 ? sw_1_0_6_down0 :
    bitdata[966:965] == 2'b10 ? cell_69_1 :
    bitdata[966:965] == 2'b01 ? cell_70_1 :
    bitdata[966:965] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[997:996] == 2'b11 ? sw_1_1_4_down0 :
    bitdata[997:996] == 2'b10 ? cell_84_0 :
    bitdata[997:996] == 2'b01 ? cell_85_0 :
    bitdata[997:996] == 2'b0 ? 8'b0 : 8'bx);
assign cell_77_0 =
   (bitdata[968:967] == 2'b11 ? sw_1_0_6_down0 :
    bitdata[968:967] == 2'b10 ? cell_69_1 :
    bitdata[968:967] == 2'b01 ? cell_70_1 :
    bitdata[968:967] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[999:998] == 2'b11 ? sw_1_1_4_down0 :
    bitdata[999:998] == 2'b10 ? cell_84_0 :
    bitdata[999:998] == 2'b01 ? cell_85_0 :
    bitdata[999:998] == 2'b0 ? 8'b0 : 8'bx);
assign cell_77_1 =
   (bitdata[970:969] == 2'b11 ? sw_1_0_6_down0 :
    bitdata[970:969] == 2'b10 ? cell_69_1 :
    bitdata[970:969] == 2'b01 ? cell_70_1 :
    bitdata[970:969] == 2'b0 ? 8'b0 : 8'bx) |
   (bitdata[1001:1000] == 2'b11 ? sw_1_1_4_down0 :
    bitdata[1001:1000] == 2'b10 ? cell_84_0 :
    bitdata[1001:1000] == 2'b01 ? cell_85_0 :
    bitdata[1001:1000] == 2'b0 ? 8'b0 : 8'bx);
assign cell_78_0 =
   (bitdata[1085:1083] == 3'b001 ? sw_2_0_5_down0 :
    bitdata[1085:1083] == 3'b100 ? cell_67_1 :
    bitdata[1085:1083] == 3'b010 ? cell_72_3 :
    bitdata[1085:1083] == 3'b110 ? cell_77_2 :
    bitdata[1085:1083] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1150:1148] == 3'b001 ? sw_2_1_4_down0 :
    bitdata[1150:1148] == 3'b100 ? cell_71_3 :
    bitdata[1150:1148] == 3'b010 ? cell_92_0 :
    bitdata[1150:1148] == 3'b110 ? cell_93_0 :
    bitdata[1150:1148] == 3'b0 ? 16'b0 : 16'bx);
assign cell_78_1 =
   (bitdata[1088:1086] == 3'b001 ? sw_2_0_5_down0 :
    bitdata[1088:1086] == 3'b100 ? cell_67_1 :
    bitdata[1088:1086] == 3'b010 ? cell_72_3 :
    bitdata[1088:1086] == 3'b110 ? cell_77_2 :
    bitdata[1088:1086] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1153:1151] == 3'b001 ? sw_2_1_4_down0 :
    bitdata[1153:1151] == 3'b100 ? cell_71_3 :
    bitdata[1153:1151] == 3'b010 ? cell_92_0 :
    bitdata[1153:1151] == 3'b110 ? cell_93_0 :
    bitdata[1153:1151] == 3'b0 ? 16'b0 : 16'bx);
assign cell_78_2 =
   (bitdata[242:242] == 1'b1 ? sw_0_0_17_down0 :
    bitdata[242:242] == 1'b0 ? 1'b0 : 1'bx) |
   (bitdata[857:855] == 3'b010 ? sw_0_1_17_down0 :
    bitdata[857:855] == 3'b110 ? sw_0_1_17_down1 :
    bitdata[857:855] == 3'b001 ? sw_0_1_17_down2 :
    bitdata[857:855] == 3'b100 ? cell_39_0 :
    bitdata[857:855] == 3'b0 ? 1'b0 : 1'bx);
assign cell_79_0 =
   (bitdata[1066:1065] == 2'b11 ? sw_2_0_4_down0 :
    bitdata[1066:1065] == 2'b10 ? cell_61_5 :
    bitdata[1066:1065] == 2'b01 ? cell_91_0 :
    bitdata[1066:1065] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1165:1163] == 3'b101 ? sw_2_1_5_down0 :
    bitdata[1165:1163] == 3'b100 ? cell_63_6 :
    bitdata[1165:1163] == 3'b010 ? cell_63_7 :
    bitdata[1165:1163] == 3'b110 ? cell_90_0 :
    bitdata[1165:1163] == 3'b001 ? cell_91_0 :
    bitdata[1165:1163] == 3'b0 ? 16'b0 : 16'bx);
assign cell_79_1 =
   (bitdata[1068:1067] == 2'b11 ? sw_2_0_4_down0 :
    bitdata[1068:1067] == 2'b10 ? cell_61_5 :
    bitdata[1068:1067] == 2'b01 ? cell_91_0 :
    bitdata[1068:1067] == 2'b0 ? 16'b0 : 16'bx) |
   (bitdata[1168:1166] == 3'b101 ? sw_2_1_5_down0 :
    bitdata[1168:1166] == 3'b100 ? cell_63_6 :
    bitdata[1168:1166] == 3'b010 ? cell_63_7 :
    bitdata[1168:1166] == 3'b110 ? cell_90_0 :
    bitdata[1168:1166] == 3'b001 ? cell_91_0 :
    bitdata[1168:1166] == 3'b0 ? 16'b0 : 16'bx);
assign cell_79_2 =
   (bitdata[238:236] == 3'b001 ? sw_0_0_16_down0 :
    bitdata[238:236] == 3'b100 ? cell_46_0 :
    bitdata[238:236] == 3'b010 ? cell_47_0 :
    bitdata[238:236] == 3'b110 ? cell_48_0 :
    bitdata[238:236] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[860:858] == 3'b010 ? sw_0_1_17_down0 :
    bitdata[860:858] == 3'b110 ? sw_0_1_17_down1 :
    bitdata[860:858] == 3'b001 ? sw_0_1_17_down2 :
    bitdata[860:858] == 3'b100 ? cell_39_0 :
    bitdata[860:858] == 3'b0 ? 1'b0 : 1'bx);
assign cell_80_0 =
   (bitdata[145:142] == 4'b1110 ? sw_0_0_8_down0 :
    bitdata[145:142] == 4'b0001 ? sw_0_0_8_down1 :
    bitdata[145:142] == 4'b1001 ? sw_0_0_8_down2 :
    bitdata[145:142] == 4'b0101 ? sw_0_0_8_down3 :
    bitdata[145:142] == 4'b1101 ? sw_0_0_8_down4 :
    bitdata[145:142] == 4'b1000 ? cell_61_6 :
    bitdata[145:142] == 4'b0100 ? cell_61_7 :
    bitdata[145:142] == 4'b1100 ? cell_71_5 :
    bitdata[145:142] == 4'b0010 ? cell_71_6 :
    bitdata[145:142] == 4'b1010 ? cell_71_7 :
    bitdata[145:142] == 4'b0110 ? cell_71_8 :
    bitdata[145:142] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[640:636] == 5'b00001 ? sw_0_1_8_down0 :
    bitdata[640:636] == 5'b10001 ? sw_0_1_8_down1 :
    bitdata[640:636] == 5'b01001 ? sw_0_1_8_down2 :
    bitdata[640:636] == 5'b11001 ? sw_0_1_8_down3 :
    bitdata[640:636] == 5'b00101 ? sw_0_1_8_down4 :
    bitdata[640:636] == 5'b10101 ? sw_0_1_8_down5 :
    bitdata[640:636] == 5'b10000 ? cell_81_10 :
    bitdata[640:636] == 5'b01000 ? cell_81_11 :
    bitdata[640:636] == 5'b11000 ? cell_81_12 :
    bitdata[640:636] == 5'b00100 ? cell_81_13 :
    bitdata[640:636] == 5'b10100 ? cell_81_14 :
    bitdata[640:636] == 5'b01100 ? cell_81_15 :
    bitdata[640:636] == 5'b11100 ? cell_81_16 :
    bitdata[640:636] == 5'b00010 ? cell_81_17 :
    bitdata[640:636] == 5'b10010 ? cell_81_18 :
    bitdata[640:636] == 5'b01010 ? cell_81_19 :
    bitdata[640:636] == 5'b11010 ? cell_81_20 :
    bitdata[640:636] == 5'b00110 ? cell_81_21 :
    bitdata[640:636] == 5'b10110 ? cell_81_22 :
    bitdata[640:636] == 5'b01110 ? cell_81_23 :
    bitdata[640:636] == 5'b11110 ? cell_81_24 :
    bitdata[640:636] == 5'b0 ? 1'b0 : 1'bx);
assign cell_80_1 =
   (bitdata[149:146] == 4'b1110 ? sw_0_0_8_down0 :
    bitdata[149:146] == 4'b0001 ? sw_0_0_8_down1 :
    bitdata[149:146] == 4'b1001 ? sw_0_0_8_down2 :
    bitdata[149:146] == 4'b0101 ? sw_0_0_8_down3 :
    bitdata[149:146] == 4'b1101 ? sw_0_0_8_down4 :
    bitdata[149:146] == 4'b1000 ? cell_61_6 :
    bitdata[149:146] == 4'b0100 ? cell_61_7 :
    bitdata[149:146] == 4'b1100 ? cell_71_5 :
    bitdata[149:146] == 4'b0010 ? cell_71_6 :
    bitdata[149:146] == 4'b1010 ? cell_71_7 :
    bitdata[149:146] == 4'b0110 ? cell_71_8 :
    bitdata[149:146] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[645:641] == 5'b00001 ? sw_0_1_8_down0 :
    bitdata[645:641] == 5'b10001 ? sw_0_1_8_down1 :
    bitdata[645:641] == 5'b01001 ? sw_0_1_8_down2 :
    bitdata[645:641] == 5'b11001 ? sw_0_1_8_down3 :
    bitdata[645:641] == 5'b00101 ? sw_0_1_8_down4 :
    bitdata[645:641] == 5'b10101 ? sw_0_1_8_down5 :
    bitdata[645:641] == 5'b10000 ? cell_81_10 :
    bitdata[645:641] == 5'b01000 ? cell_81_11 :
    bitdata[645:641] == 5'b11000 ? cell_81_12 :
    bitdata[645:641] == 5'b00100 ? cell_81_13 :
    bitdata[645:641] == 5'b10100 ? cell_81_14 :
    bitdata[645:641] == 5'b01100 ? cell_81_15 :
    bitdata[645:641] == 5'b11100 ? cell_81_16 :
    bitdata[645:641] == 5'b00010 ? cell_81_17 :
    bitdata[645:641] == 5'b10010 ? cell_81_18 :
    bitdata[645:641] == 5'b01010 ? cell_81_19 :
    bitdata[645:641] == 5'b11010 ? cell_81_20 :
    bitdata[645:641] == 5'b00110 ? cell_81_21 :
    bitdata[645:641] == 5'b10110 ? cell_81_22 :
    bitdata[645:641] == 5'b01110 ? cell_81_23 :
    bitdata[645:641] == 5'b11110 ? cell_81_24 :
    bitdata[645:641] == 5'b0 ? 1'b0 : 1'bx);
assign cell_80_2 =
   (bitdata[153:150] == 4'b1110 ? sw_0_0_8_down0 :
    bitdata[153:150] == 4'b0001 ? sw_0_0_8_down1 :
    bitdata[153:150] == 4'b1001 ? sw_0_0_8_down2 :
    bitdata[153:150] == 4'b0101 ? sw_0_0_8_down3 :
    bitdata[153:150] == 4'b1101 ? sw_0_0_8_down4 :
    bitdata[153:150] == 4'b1000 ? cell_61_6 :
    bitdata[153:150] == 4'b0100 ? cell_61_7 :
    bitdata[153:150] == 4'b1100 ? cell_71_5 :
    bitdata[153:150] == 4'b0010 ? cell_71_6 :
    bitdata[153:150] == 4'b1010 ? cell_71_7 :
    bitdata[153:150] == 4'b0110 ? cell_71_8 :
    bitdata[153:150] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[650:646] == 5'b00001 ? sw_0_1_8_down0 :
    bitdata[650:646] == 5'b10001 ? sw_0_1_8_down1 :
    bitdata[650:646] == 5'b01001 ? sw_0_1_8_down2 :
    bitdata[650:646] == 5'b11001 ? sw_0_1_8_down3 :
    bitdata[650:646] == 5'b00101 ? sw_0_1_8_down4 :
    bitdata[650:646] == 5'b10101 ? sw_0_1_8_down5 :
    bitdata[650:646] == 5'b10000 ? cell_81_10 :
    bitdata[650:646] == 5'b01000 ? cell_81_11 :
    bitdata[650:646] == 5'b11000 ? cell_81_12 :
    bitdata[650:646] == 5'b00100 ? cell_81_13 :
    bitdata[650:646] == 5'b10100 ? cell_81_14 :
    bitdata[650:646] == 5'b01100 ? cell_81_15 :
    bitdata[650:646] == 5'b11100 ? cell_81_16 :
    bitdata[650:646] == 5'b00010 ? cell_81_17 :
    bitdata[650:646] == 5'b10010 ? cell_81_18 :
    bitdata[650:646] == 5'b01010 ? cell_81_19 :
    bitdata[650:646] == 5'b11010 ? cell_81_20 :
    bitdata[650:646] == 5'b00110 ? cell_81_21 :
    bitdata[650:646] == 5'b10110 ? cell_81_22 :
    bitdata[650:646] == 5'b01110 ? cell_81_23 :
    bitdata[650:646] == 5'b11110 ? cell_81_24 :
    bitdata[650:646] == 5'b0 ? 1'b0 : 1'bx);
assign cell_80_3 =
   (bitdata[157:154] == 4'b1110 ? sw_0_0_8_down0 :
    bitdata[157:154] == 4'b0001 ? sw_0_0_8_down1 :
    bitdata[157:154] == 4'b1001 ? sw_0_0_8_down2 :
    bitdata[157:154] == 4'b0101 ? sw_0_0_8_down3 :
    bitdata[157:154] == 4'b1101 ? sw_0_0_8_down4 :
    bitdata[157:154] == 4'b1000 ? cell_61_6 :
    bitdata[157:154] == 4'b0100 ? cell_61_7 :
    bitdata[157:154] == 4'b1100 ? cell_71_5 :
    bitdata[157:154] == 4'b0010 ? cell_71_6 :
    bitdata[157:154] == 4'b1010 ? cell_71_7 :
    bitdata[157:154] == 4'b0110 ? cell_71_8 :
    bitdata[157:154] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[655:651] == 5'b00001 ? sw_0_1_8_down0 :
    bitdata[655:651] == 5'b10001 ? sw_0_1_8_down1 :
    bitdata[655:651] == 5'b01001 ? sw_0_1_8_down2 :
    bitdata[655:651] == 5'b11001 ? sw_0_1_8_down3 :
    bitdata[655:651] == 5'b00101 ? sw_0_1_8_down4 :
    bitdata[655:651] == 5'b10101 ? sw_0_1_8_down5 :
    bitdata[655:651] == 5'b10000 ? cell_81_10 :
    bitdata[655:651] == 5'b01000 ? cell_81_11 :
    bitdata[655:651] == 5'b11000 ? cell_81_12 :
    bitdata[655:651] == 5'b00100 ? cell_81_13 :
    bitdata[655:651] == 5'b10100 ? cell_81_14 :
    bitdata[655:651] == 5'b01100 ? cell_81_15 :
    bitdata[655:651] == 5'b11100 ? cell_81_16 :
    bitdata[655:651] == 5'b00010 ? cell_81_17 :
    bitdata[655:651] == 5'b10010 ? cell_81_18 :
    bitdata[655:651] == 5'b01010 ? cell_81_19 :
    bitdata[655:651] == 5'b11010 ? cell_81_20 :
    bitdata[655:651] == 5'b00110 ? cell_81_21 :
    bitdata[655:651] == 5'b10110 ? cell_81_22 :
    bitdata[655:651] == 5'b01110 ? cell_81_23 :
    bitdata[655:651] == 5'b11110 ? cell_81_24 :
    bitdata[655:651] == 5'b0 ? 1'b0 : 1'bx);
assign cell_80_4 =
   (bitdata[161:158] == 4'b1110 ? sw_0_0_8_down0 :
    bitdata[161:158] == 4'b0001 ? sw_0_0_8_down1 :
    bitdata[161:158] == 4'b1001 ? sw_0_0_8_down2 :
    bitdata[161:158] == 4'b0101 ? sw_0_0_8_down3 :
    bitdata[161:158] == 4'b1101 ? sw_0_0_8_down4 :
    bitdata[161:158] == 4'b1000 ? cell_61_6 :
    bitdata[161:158] == 4'b0100 ? cell_61_7 :
    bitdata[161:158] == 4'b1100 ? cell_71_5 :
    bitdata[161:158] == 4'b0010 ? cell_71_6 :
    bitdata[161:158] == 4'b1010 ? cell_71_7 :
    bitdata[161:158] == 4'b0110 ? cell_71_8 :
    bitdata[161:158] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[660:656] == 5'b00001 ? sw_0_1_8_down0 :
    bitdata[660:656] == 5'b10001 ? sw_0_1_8_down1 :
    bitdata[660:656] == 5'b01001 ? sw_0_1_8_down2 :
    bitdata[660:656] == 5'b11001 ? sw_0_1_8_down3 :
    bitdata[660:656] == 5'b00101 ? sw_0_1_8_down4 :
    bitdata[660:656] == 5'b10101 ? sw_0_1_8_down5 :
    bitdata[660:656] == 5'b10000 ? cell_81_10 :
    bitdata[660:656] == 5'b01000 ? cell_81_11 :
    bitdata[660:656] == 5'b11000 ? cell_81_12 :
    bitdata[660:656] == 5'b00100 ? cell_81_13 :
    bitdata[660:656] == 5'b10100 ? cell_81_14 :
    bitdata[660:656] == 5'b01100 ? cell_81_15 :
    bitdata[660:656] == 5'b11100 ? cell_81_16 :
    bitdata[660:656] == 5'b00010 ? cell_81_17 :
    bitdata[660:656] == 5'b10010 ? cell_81_18 :
    bitdata[660:656] == 5'b01010 ? cell_81_19 :
    bitdata[660:656] == 5'b11010 ? cell_81_20 :
    bitdata[660:656] == 5'b00110 ? cell_81_21 :
    bitdata[660:656] == 5'b10110 ? cell_81_22 :
    bitdata[660:656] == 5'b01110 ? cell_81_23 :
    bitdata[660:656] == 5'b11110 ? cell_81_24 :
    bitdata[660:656] == 5'b0 ? 1'b0 : 1'bx);
assign cell_80_5 =
   (bitdata[165:162] == 4'b1110 ? sw_0_0_8_down0 :
    bitdata[165:162] == 4'b0001 ? sw_0_0_8_down1 :
    bitdata[165:162] == 4'b1001 ? sw_0_0_8_down2 :
    bitdata[165:162] == 4'b0101 ? sw_0_0_8_down3 :
    bitdata[165:162] == 4'b1101 ? sw_0_0_8_down4 :
    bitdata[165:162] == 4'b1000 ? cell_61_6 :
    bitdata[165:162] == 4'b0100 ? cell_61_7 :
    bitdata[165:162] == 4'b1100 ? cell_71_5 :
    bitdata[165:162] == 4'b0010 ? cell_71_6 :
    bitdata[165:162] == 4'b1010 ? cell_71_7 :
    bitdata[165:162] == 4'b0110 ? cell_71_8 :
    bitdata[165:162] == 4'b0 ? 1'b0 : 1'bx) |
   (bitdata[665:661] == 5'b00001 ? sw_0_1_8_down0 :
    bitdata[665:661] == 5'b10001 ? sw_0_1_8_down1 :
    bitdata[665:661] == 5'b01001 ? sw_0_1_8_down2 :
    bitdata[665:661] == 5'b11001 ? sw_0_1_8_down3 :
    bitdata[665:661] == 5'b00101 ? sw_0_1_8_down4 :
    bitdata[665:661] == 5'b10101 ? sw_0_1_8_down5 :
    bitdata[665:661] == 5'b10000 ? cell_81_10 :
    bitdata[665:661] == 5'b01000 ? cell_81_11 :
    bitdata[665:661] == 5'b11000 ? cell_81_12 :
    bitdata[665:661] == 5'b00100 ? cell_81_13 :
    bitdata[665:661] == 5'b10100 ? cell_81_14 :
    bitdata[665:661] == 5'b01100 ? cell_81_15 :
    bitdata[665:661] == 5'b11100 ? cell_81_16 :
    bitdata[665:661] == 5'b00010 ? cell_81_17 :
    bitdata[665:661] == 5'b10010 ? cell_81_18 :
    bitdata[665:661] == 5'b01010 ? cell_81_19 :
    bitdata[665:661] == 5'b11010 ? cell_81_20 :
    bitdata[665:661] == 5'b00110 ? cell_81_21 :
    bitdata[665:661] == 5'b10110 ? cell_81_22 :
    bitdata[665:661] == 5'b01110 ? cell_81_23 :
    bitdata[665:661] == 5'b11110 ? cell_81_24 :
    bitdata[665:661] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_0 =
   (bitdata[340:338] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[340:338] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[340:338] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[340:338] == 3'b100 ? cell_63_8 :
    bitdata[340:338] == 3'b010 ? cell_63_9 :
    bitdata[340:338] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[670:666] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[670:666] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[670:666] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[670:666] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[670:666] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[670:666] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[670:666] == 5'b10000 ? cell_80_6 :
    bitdata[670:666] == 5'b01000 ? cell_80_7 :
    bitdata[670:666] == 5'b11000 ? cell_80_8 :
    bitdata[670:666] == 5'b00100 ? cell_80_9 :
    bitdata[670:666] == 5'b10100 ? cell_80_10 :
    bitdata[670:666] == 5'b01100 ? cell_80_11 :
    bitdata[670:666] == 5'b11100 ? cell_80_12 :
    bitdata[670:666] == 5'b00010 ? cell_80_13 :
    bitdata[670:666] == 5'b10010 ? cell_80_14 :
    bitdata[670:666] == 5'b01010 ? cell_80_15 :
    bitdata[670:666] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_1 =
   (bitdata[343:341] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[343:341] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[343:341] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[343:341] == 3'b100 ? cell_63_8 :
    bitdata[343:341] == 3'b010 ? cell_63_9 :
    bitdata[343:341] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[675:671] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[675:671] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[675:671] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[675:671] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[675:671] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[675:671] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[675:671] == 5'b10000 ? cell_80_6 :
    bitdata[675:671] == 5'b01000 ? cell_80_7 :
    bitdata[675:671] == 5'b11000 ? cell_80_8 :
    bitdata[675:671] == 5'b00100 ? cell_80_9 :
    bitdata[675:671] == 5'b10100 ? cell_80_10 :
    bitdata[675:671] == 5'b01100 ? cell_80_11 :
    bitdata[675:671] == 5'b11100 ? cell_80_12 :
    bitdata[675:671] == 5'b00010 ? cell_80_13 :
    bitdata[675:671] == 5'b10010 ? cell_80_14 :
    bitdata[675:671] == 5'b01010 ? cell_80_15 :
    bitdata[675:671] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_2 =
   (bitdata[346:344] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[346:344] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[346:344] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[346:344] == 3'b100 ? cell_63_8 :
    bitdata[346:344] == 3'b010 ? cell_63_9 :
    bitdata[346:344] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[680:676] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[680:676] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[680:676] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[680:676] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[680:676] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[680:676] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[680:676] == 5'b10000 ? cell_80_6 :
    bitdata[680:676] == 5'b01000 ? cell_80_7 :
    bitdata[680:676] == 5'b11000 ? cell_80_8 :
    bitdata[680:676] == 5'b00100 ? cell_80_9 :
    bitdata[680:676] == 5'b10100 ? cell_80_10 :
    bitdata[680:676] == 5'b01100 ? cell_80_11 :
    bitdata[680:676] == 5'b11100 ? cell_80_12 :
    bitdata[680:676] == 5'b00010 ? cell_80_13 :
    bitdata[680:676] == 5'b10010 ? cell_80_14 :
    bitdata[680:676] == 5'b01010 ? cell_80_15 :
    bitdata[680:676] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_3 =
   (bitdata[349:347] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[349:347] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[349:347] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[349:347] == 3'b100 ? cell_63_8 :
    bitdata[349:347] == 3'b010 ? cell_63_9 :
    bitdata[349:347] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[685:681] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[685:681] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[685:681] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[685:681] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[685:681] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[685:681] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[685:681] == 5'b10000 ? cell_80_6 :
    bitdata[685:681] == 5'b01000 ? cell_80_7 :
    bitdata[685:681] == 5'b11000 ? cell_80_8 :
    bitdata[685:681] == 5'b00100 ? cell_80_9 :
    bitdata[685:681] == 5'b10100 ? cell_80_10 :
    bitdata[685:681] == 5'b01100 ? cell_80_11 :
    bitdata[685:681] == 5'b11100 ? cell_80_12 :
    bitdata[685:681] == 5'b00010 ? cell_80_13 :
    bitdata[685:681] == 5'b10010 ? cell_80_14 :
    bitdata[685:681] == 5'b01010 ? cell_80_15 :
    bitdata[685:681] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_4 =
   (bitdata[352:350] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[352:350] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[352:350] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[352:350] == 3'b100 ? cell_63_8 :
    bitdata[352:350] == 3'b010 ? cell_63_9 :
    bitdata[352:350] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[690:686] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[690:686] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[690:686] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[690:686] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[690:686] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[690:686] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[690:686] == 5'b10000 ? cell_80_6 :
    bitdata[690:686] == 5'b01000 ? cell_80_7 :
    bitdata[690:686] == 5'b11000 ? cell_80_8 :
    bitdata[690:686] == 5'b00100 ? cell_80_9 :
    bitdata[690:686] == 5'b10100 ? cell_80_10 :
    bitdata[690:686] == 5'b01100 ? cell_80_11 :
    bitdata[690:686] == 5'b11100 ? cell_80_12 :
    bitdata[690:686] == 5'b00010 ? cell_80_13 :
    bitdata[690:686] == 5'b10010 ? cell_80_14 :
    bitdata[690:686] == 5'b01010 ? cell_80_15 :
    bitdata[690:686] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_5 =
   (bitdata[355:353] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[355:353] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[355:353] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[355:353] == 3'b100 ? cell_63_8 :
    bitdata[355:353] == 3'b010 ? cell_63_9 :
    bitdata[355:353] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[695:691] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[695:691] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[695:691] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[695:691] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[695:691] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[695:691] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[695:691] == 5'b10000 ? cell_80_6 :
    bitdata[695:691] == 5'b01000 ? cell_80_7 :
    bitdata[695:691] == 5'b11000 ? cell_80_8 :
    bitdata[695:691] == 5'b00100 ? cell_80_9 :
    bitdata[695:691] == 5'b10100 ? cell_80_10 :
    bitdata[695:691] == 5'b01100 ? cell_80_11 :
    bitdata[695:691] == 5'b11100 ? cell_80_12 :
    bitdata[695:691] == 5'b00010 ? cell_80_13 :
    bitdata[695:691] == 5'b10010 ? cell_80_14 :
    bitdata[695:691] == 5'b01010 ? cell_80_15 :
    bitdata[695:691] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_6 =
   (bitdata[358:356] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[358:356] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[358:356] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[358:356] == 3'b100 ? cell_63_8 :
    bitdata[358:356] == 3'b010 ? cell_63_9 :
    bitdata[358:356] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[700:696] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[700:696] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[700:696] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[700:696] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[700:696] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[700:696] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[700:696] == 5'b10000 ? cell_80_6 :
    bitdata[700:696] == 5'b01000 ? cell_80_7 :
    bitdata[700:696] == 5'b11000 ? cell_80_8 :
    bitdata[700:696] == 5'b00100 ? cell_80_9 :
    bitdata[700:696] == 5'b10100 ? cell_80_10 :
    bitdata[700:696] == 5'b01100 ? cell_80_11 :
    bitdata[700:696] == 5'b11100 ? cell_80_12 :
    bitdata[700:696] == 5'b00010 ? cell_80_13 :
    bitdata[700:696] == 5'b10010 ? cell_80_14 :
    bitdata[700:696] == 5'b01010 ? cell_80_15 :
    bitdata[700:696] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_7 =
   (bitdata[361:359] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[361:359] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[361:359] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[361:359] == 3'b100 ? cell_63_8 :
    bitdata[361:359] == 3'b010 ? cell_63_9 :
    bitdata[361:359] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[705:701] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[705:701] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[705:701] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[705:701] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[705:701] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[705:701] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[705:701] == 5'b10000 ? cell_80_6 :
    bitdata[705:701] == 5'b01000 ? cell_80_7 :
    bitdata[705:701] == 5'b11000 ? cell_80_8 :
    bitdata[705:701] == 5'b00100 ? cell_80_9 :
    bitdata[705:701] == 5'b10100 ? cell_80_10 :
    bitdata[705:701] == 5'b01100 ? cell_80_11 :
    bitdata[705:701] == 5'b11100 ? cell_80_12 :
    bitdata[705:701] == 5'b00010 ? cell_80_13 :
    bitdata[705:701] == 5'b10010 ? cell_80_14 :
    bitdata[705:701] == 5'b01010 ? cell_80_15 :
    bitdata[705:701] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_8 =
   (bitdata[364:362] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[364:362] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[364:362] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[364:362] == 3'b100 ? cell_63_8 :
    bitdata[364:362] == 3'b010 ? cell_63_9 :
    bitdata[364:362] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[710:706] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[710:706] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[710:706] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[710:706] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[710:706] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[710:706] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[710:706] == 5'b10000 ? cell_80_6 :
    bitdata[710:706] == 5'b01000 ? cell_80_7 :
    bitdata[710:706] == 5'b11000 ? cell_80_8 :
    bitdata[710:706] == 5'b00100 ? cell_80_9 :
    bitdata[710:706] == 5'b10100 ? cell_80_10 :
    bitdata[710:706] == 5'b01100 ? cell_80_11 :
    bitdata[710:706] == 5'b11100 ? cell_80_12 :
    bitdata[710:706] == 5'b00010 ? cell_80_13 :
    bitdata[710:706] == 5'b10010 ? cell_80_14 :
    bitdata[710:706] == 5'b01010 ? cell_80_15 :
    bitdata[710:706] == 5'b0 ? 1'b0 : 1'bx);
assign cell_81_9 =
   (bitdata[367:365] == 3'b110 ? sw_0_0_25_down0 :
    bitdata[367:365] == 3'b001 ? sw_0_0_25_down1 :
    bitdata[367:365] == 3'b101 ? sw_0_0_25_down2 :
    bitdata[367:365] == 3'b100 ? cell_63_8 :
    bitdata[367:365] == 3'b010 ? cell_63_9 :
    bitdata[367:365] == 3'b0 ? 1'b0 : 1'bx) |
   (bitdata[715:711] == 5'b11010 ? sw_0_1_8_down0 :
    bitdata[715:711] == 5'b00110 ? sw_0_1_8_down1 :
    bitdata[715:711] == 5'b10110 ? sw_0_1_8_down2 :
    bitdata[715:711] == 5'b01110 ? sw_0_1_8_down3 :
    bitdata[715:711] == 5'b11110 ? sw_0_1_8_down4 :
    bitdata[715:711] == 5'b00001 ? sw_0_1_8_down5 :
    bitdata[715:711] == 5'b10000 ? cell_80_6 :
    bitdata[715:711] == 5'b01000 ? cell_80_7 :
    bitdata[715:711] == 5'b11000 ? cell_80_8 :
    bitdata[715:711] == 5'b00100 ? cell_80_9 :
    bitdata[715:711] == 5'b10100 ? cell_80_10 :
    bitdata[715:711] == 5'b01100 ? cell_80_11 :
    bitdata[715:711] == 5'b11100 ? cell_80_12 :
    bitdata[715:711] == 5'b00010 ? cell_80_13 :
    bitdata[715:711] == 5'b10010 ? cell_80_14 :
    bitdata[715:711] == 5'b01010 ? cell_80_15 :
    bitdata[715:711] == 5'b0 ? 1'b0 : 1'bx);
assign cell_96_0 =
   (bitdata[1112:1110] == 3'b001 ? sw_2_0_7_down0 :
    bitdata[1112:1110] == 3'b100 ? cell_65_2 :
    bitdata[1112:1110] == 3'b010 ? cell_66_1 :
    bitdata[1112:1110] == 3'b110 ? cell_71_3 :
    bitdata[1112:1110] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1137:1136] == 2'b11 ? sw_2_1_3_down0 :
    bitdata[1137:1136] == 2'b10 ? cell_94_0 :
    bitdata[1137:1136] == 2'b01 ? cell_95_0 :
    bitdata[1137:1136] == 2'b0 ? 16'b0 : 16'bx);
assign cell_97_0 =
   (bitdata[1071:1069] == 3'b001 ? sw_2_0_4_down0 :
    bitdata[1071:1069] == 3'b100 ? cell_61_5 :
    bitdata[1071:1069] == 3'b010 ? cell_79_3 :
    bitdata[1071:1069] == 3'b110 ? cell_91_0 :
    bitdata[1071:1069] == 3'b0 ? 16'b0 : 16'bx) |
   (bitdata[1139:1138] == 2'b11 ? sw_2_1_3_down0 :
    bitdata[1139:1138] == 2'b10 ? cell_94_0 :
    bitdata[1139:1138] == 2'b01 ? cell_95_0 :
    bitdata[1139:1138] == 2'b0 ? 16'b0 : 16'bx);
assign cell_9_0 =
   (bitdata[302:298] == 5'b01001 ? sw_0_0_25_down0 :
    bitdata[302:298] == 5'b11001 ? sw_0_0_25_down1 :
    bitdata[302:298] == 5'b00101 ? sw_0_0_25_down2 :
    bitdata[302:298] == 5'b10000 ? cell_63_8 :
    bitdata[302:298] == 5'b01000 ? cell_63_9 :
    bitdata[302:298] == 5'b11000 ? cell_81_10 :
    bitdata[302:298] == 5'b00100 ? cell_81_11 :
    bitdata[302:298] == 5'b10100 ? cell_81_12 :
    bitdata[302:298] == 5'b01100 ? cell_81_13 :
    bitdata[302:298] == 5'b11100 ? cell_81_14 :
    bitdata[302:298] == 5'b00010 ? cell_81_15 :
    bitdata[302:298] == 5'b10010 ? cell_81_16 :
    bitdata[302:298] == 5'b01010 ? cell_81_17 :
    bitdata[302:298] == 5'b11010 ? cell_81_18 :
    bitdata[302:298] == 5'b00110 ? cell_81_19 :
    bitdata[302:298] == 5'b10110 ? cell_81_20 :
    bitdata[302:298] == 5'b01110 ? cell_81_21 :
    bitdata[302:298] == 5'b11110 ? cell_81_22 :
    bitdata[302:298] == 5'b00001 ? cell_81_23 :
    bitdata[302:298] == 5'b10001 ? cell_81_24 :
    bitdata[302:298] == 5'b0 ? 1'b0 : 1'bx) |
   (bitdata[907:905] == 3'b001 ? sw_0_1_25_down0 :
    bitdata[907:905] == 3'b100 ? cell_6_0 :
    bitdata[907:905] == 3'b010 ? cell_7_0 :
    bitdata[907:905] == 3'b110 ? cell_8_0 :
    bitdata[907:905] == 3'b0 ? 1'b0 : 1'bx);
assign sw_0_0_10_down0 =
   (bitdata[33:30] == 4'b0001 ? sw_0_0_3_down0 :
    bitdata[33:30] == 4'b0000 ? sw_0_0_8_up0 :
    bitdata[33:30] == 4'b1000 ? sw_0_0_8_up1 :
    bitdata[33:30] == 4'b0100 ? sw_0_0_8_up2 :
    bitdata[33:30] == 4'b1100 ? sw_0_0_9_up0 :
    bitdata[33:30] == 4'b0010 ? sw_0_0_9_up1 :
    bitdata[33:30] == 4'b1010 ? sw_0_0_9_up2 :
    bitdata[33:30] == 4'b0110 ? sw_0_0_9_up3 :
    bitdata[33:30] == 4'b1110 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_10_down1 =
   (bitdata[37:34] == 4'b0001 ? sw_0_0_3_down0 :
    bitdata[37:34] == 4'b0000 ? sw_0_0_8_up0 :
    bitdata[37:34] == 4'b1000 ? sw_0_0_8_up1 :
    bitdata[37:34] == 4'b0100 ? sw_0_0_8_up2 :
    bitdata[37:34] == 4'b1100 ? sw_0_0_9_up0 :
    bitdata[37:34] == 4'b0010 ? sw_0_0_9_up1 :
    bitdata[37:34] == 4'b1010 ? sw_0_0_9_up2 :
    bitdata[37:34] == 4'b0110 ? sw_0_0_9_up3 :
    bitdata[37:34] == 4'b1110 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_10_down2 =
   (bitdata[41:38] == 4'b0001 ? sw_0_0_3_down0 :
    bitdata[41:38] == 4'b0000 ? sw_0_0_8_up0 :
    bitdata[41:38] == 4'b1000 ? sw_0_0_8_up1 :
    bitdata[41:38] == 4'b0100 ? sw_0_0_8_up2 :
    bitdata[41:38] == 4'b1100 ? sw_0_0_9_up0 :
    bitdata[41:38] == 4'b0010 ? sw_0_0_9_up1 :
    bitdata[41:38] == 4'b1010 ? sw_0_0_9_up2 :
    bitdata[41:38] == 4'b0110 ? sw_0_0_9_up3 :
    bitdata[41:38] == 4'b1110 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_10_up0 =
   (bitdata[176:174] == 3'b000 ? cell_62_6 :
    bitdata[176:174] == 3'b100 ? cell_62_7 :
    bitdata[176:174] == 3'b010 ? cell_64_8 :
    bitdata[176:174] == 3'b110 ? cell_64_9 :
    bitdata[176:174] == 3'b001 ? cell_83_0 : 1'bx);
assign sw_0_0_11_down0 =
   (bitdata[45:42] == 4'b0001 ? sw_0_0_3_down0 :
    bitdata[45:42] == 4'b0000 ? sw_0_0_8_up0 :
    bitdata[45:42] == 4'b1000 ? sw_0_0_8_up1 :
    bitdata[45:42] == 4'b0100 ? sw_0_0_8_up2 :
    bitdata[45:42] == 4'b1100 ? sw_0_0_9_up0 :
    bitdata[45:42] == 4'b0010 ? sw_0_0_9_up1 :
    bitdata[45:42] == 4'b1010 ? sw_0_0_9_up2 :
    bitdata[45:42] == 4'b0110 ? sw_0_0_9_up3 :
    bitdata[45:42] == 4'b1110 ? sw_0_0_10_up0 : 1'bx);
assign sw_0_0_11_down1 =
   (bitdata[49:46] == 4'b0001 ? sw_0_0_3_down0 :
    bitdata[49:46] == 4'b0000 ? sw_0_0_8_up0 :
    bitdata[49:46] == 4'b1000 ? sw_0_0_8_up1 :
    bitdata[49:46] == 4'b0100 ? sw_0_0_8_up2 :
    bitdata[49:46] == 4'b1100 ? sw_0_0_9_up0 :
    bitdata[49:46] == 4'b0010 ? sw_0_0_9_up1 :
    bitdata[49:46] == 4'b1010 ? sw_0_0_9_up2 :
    bitdata[49:46] == 4'b0110 ? sw_0_0_9_up3 :
    bitdata[49:46] == 4'b1110 ? sw_0_0_10_up0 : 1'bx);
assign sw_0_0_11_up0 = cell_43_0;
assign sw_0_0_12_down0 =
   (bitdata[51:51] == 1'b1 ? sw_0_0_4_down0 :
    bitdata[51:51] == 1'b0 ? sw_0_0_15_up0 : 1'bx);
assign sw_0_0_12_up0 =
   (bitdata[213:211] == 3'b000 ? cell_8_0 :
    bitdata[213:211] == 3'b100 ? cell_72_5 :
    bitdata[213:211] == 3'b010 ? cell_72_6 :
    bitdata[213:211] == 3'b110 ? cell_72_7 :
    bitdata[213:211] == 3'b001 ? cell_72_8 : 1'bx);
assign sw_0_0_13_down0 =
   (bitdata[53:52] == 2'b01 ? sw_0_0_4_down0 :
    bitdata[53:52] == 2'b00 ? sw_0_0_12_up0 :
    bitdata[53:52] == 2'b10 ? sw_0_0_15_up0 : 1'bx);
assign sw_0_0_14_down0 =
   (bitdata[55:54] == 2'b01 ? sw_0_0_4_down0 :
    bitdata[55:54] == 2'b00 ? sw_0_0_12_up0 :
    bitdata[55:54] == 2'b10 ? sw_0_0_15_up0 : 1'bx);
assign sw_0_0_15_up0 =
   (bitdata[233:232] == 2'b00 ? cell_49_0 :
    bitdata[233:232] == 2'b10 ? cell_50_0 :
    bitdata[233:232] == 2'b01 ? cell_51_0 :
    bitdata[233:232] == 2'b11 ? cell_52_0 : 1'bx);
assign sw_0_0_16_down0 =
   (bitdata[57:57] == 1'b1 ? sw_0_0_5_down0 :
    bitdata[57:57] == 1'b0 ? sw_0_0_18_up0 : 1'bx);
assign sw_0_0_16_up0 =
   (bitdata[235:234] == 2'b00 ? cell_46_0 :
    bitdata[235:234] == 2'b10 ? cell_47_0 :
    bitdata[235:234] == 2'b01 ? cell_48_0 : 1'bx);
assign sw_0_0_17_down0 =
   (bitdata[59:58] == 2'b01 ? sw_0_0_5_down0 :
    bitdata[59:58] == 2'b00 ? sw_0_0_16_up0 :
    bitdata[59:58] == 2'b10 ? sw_0_0_18_up0 : 1'bx);
assign sw_0_0_18_down0 =
   (bitdata[60:60] == 1'b1 ? sw_0_0_5_down0 :
    bitdata[60:60] == 1'b0 ? sw_0_0_16_up0 : 1'bx);
assign sw_0_0_18_up0 =
   (bitdata[243:243] == 1'b0 ? cell_39_0 :
    bitdata[243:243] == 1'b1 ? cell_40_0 : 1'bx);
assign sw_0_0_19_down0 =
   (bitdata[62:61] == 2'b01 ? sw_0_0_5_down0 :
    bitdata[62:61] == 2'b00 ? sw_0_0_16_up0 :
    bitdata[62:61] == 2'b10 ? sw_0_0_18_up0 : 1'bx);
assign sw_0_0_1_down0 = sw_0_0_2_up0;
assign sw_0_0_1_up0 =
   (bitdata[1:0] == 2'b00 ? sw_0_0_3_up0 :
    bitdata[1:0] == 2'b10 ? sw_0_0_4_up0 :
    bitdata[1:0] == 2'b01 ? sw_0_0_5_up0 : 1'bx);
assign sw_0_0_20_down0 =
   (bitdata[66:65] == 2'b01 ? sw_0_0_6_down0 :
    bitdata[66:65] == 2'b00 ? sw_0_0_22_up0 :
    bitdata[66:65] == 2'b10 ? sw_0_0_23_up0 : 1'bx);
assign sw_0_0_20_up0 = cell_7_0;
assign sw_0_0_21_down0 =
   (bitdata[68:67] == 2'b11 ? sw_0_0_6_down0 :
    bitdata[68:67] == 2'b00 ? sw_0_0_20_up0 :
    bitdata[68:67] == 2'b10 ? sw_0_0_22_up0 :
    bitdata[68:67] == 2'b01 ? sw_0_0_23_up0 : 1'bx);
assign sw_0_0_22_down0 =
   (bitdata[70:69] == 2'b01 ? sw_0_0_6_down0 :
    bitdata[70:69] == 2'b00 ? sw_0_0_20_up0 :
    bitdata[70:69] == 2'b10 ? sw_0_0_23_up0 : 1'bx);
assign sw_0_0_22_up0 =
   (bitdata[263:262] == 2'b00 ? cell_19_0 :
    bitdata[263:262] == 2'b10 ? cell_20_0 :
    bitdata[263:262] == 2'b01 ? cell_21_0 : 1'bx);
assign sw_0_0_23_up0 =
   (bitdata[268:267] == 2'b00 ? cell_15_0 :
    bitdata[268:267] == 2'b10 ? cell_16_0 :
    bitdata[268:267] == 2'b01 ? cell_17_0 :
    bitdata[268:267] == 2'b11 ? cell_18_0 : 1'bx);
assign sw_0_0_24_down0 =
   (bitdata[76:74] == 3'b101 ? sw_0_0_7_down0 :
    bitdata[76:74] == 3'b000 ? sw_0_0_25_up0 :
    bitdata[76:74] == 3'b100 ? sw_0_0_25_up1 :
    bitdata[76:74] == 3'b010 ? sw_0_0_25_up2 :
    bitdata[76:74] == 3'b110 ? sw_0_0_25_up3 :
    bitdata[76:74] == 3'b001 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_24_down1 =
   (bitdata[79:77] == 3'b101 ? sw_0_0_7_down0 :
    bitdata[79:77] == 3'b000 ? sw_0_0_25_up0 :
    bitdata[79:77] == 3'b100 ? sw_0_0_25_up1 :
    bitdata[79:77] == 3'b010 ? sw_0_0_25_up2 :
    bitdata[79:77] == 3'b110 ? sw_0_0_25_up3 :
    bitdata[79:77] == 3'b001 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_24_down2 =
   (bitdata[82:80] == 3'b101 ? sw_0_0_7_down0 :
    bitdata[82:80] == 3'b000 ? sw_0_0_25_up0 :
    bitdata[82:80] == 3'b100 ? sw_0_0_25_up1 :
    bitdata[82:80] == 3'b010 ? sw_0_0_25_up2 :
    bitdata[82:80] == 3'b110 ? sw_0_0_25_up3 :
    bitdata[82:80] == 3'b001 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_24_up0 = cell_3_0;
assign sw_0_0_25_down0 =
   (bitdata[84:83] == 2'b01 ? sw_0_0_7_down0 :
    bitdata[84:83] == 2'b00 ? sw_0_0_24_up0 :
    bitdata[84:83] == 2'b10 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_25_down1 =
   (bitdata[86:85] == 2'b01 ? sw_0_0_7_down0 :
    bitdata[86:85] == 2'b00 ? sw_0_0_24_up0 :
    bitdata[86:85] == 2'b10 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_25_down2 =
   (bitdata[88:87] == 2'b01 ? sw_0_0_7_down0 :
    bitdata[88:87] == 2'b00 ? sw_0_0_24_up0 :
    bitdata[88:87] == 2'b10 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_25_up0 =
   (bitdata[282:278] == 5'b00000 ? cell_63_8 :
    bitdata[282:278] == 5'b10000 ? cell_63_9 :
    bitdata[282:278] == 5'b01000 ? cell_81_10 :
    bitdata[282:278] == 5'b11000 ? cell_81_11 :
    bitdata[282:278] == 5'b00100 ? cell_81_12 :
    bitdata[282:278] == 5'b10100 ? cell_81_13 :
    bitdata[282:278] == 5'b01100 ? cell_81_14 :
    bitdata[282:278] == 5'b11100 ? cell_81_15 :
    bitdata[282:278] == 5'b00010 ? cell_81_16 :
    bitdata[282:278] == 5'b10010 ? cell_81_17 :
    bitdata[282:278] == 5'b01010 ? cell_81_18 :
    bitdata[282:278] == 5'b11010 ? cell_81_19 :
    bitdata[282:278] == 5'b00110 ? cell_81_20 :
    bitdata[282:278] == 5'b10110 ? cell_81_21 :
    bitdata[282:278] == 5'b01110 ? cell_81_22 :
    bitdata[282:278] == 5'b11110 ? cell_81_23 :
    bitdata[282:278] == 5'b00001 ? cell_81_24 : 1'bx);
assign sw_0_0_25_up1 =
   (bitdata[287:283] == 5'b00000 ? cell_63_8 :
    bitdata[287:283] == 5'b10000 ? cell_63_9 :
    bitdata[287:283] == 5'b01000 ? cell_81_10 :
    bitdata[287:283] == 5'b11000 ? cell_81_11 :
    bitdata[287:283] == 5'b00100 ? cell_81_12 :
    bitdata[287:283] == 5'b10100 ? cell_81_13 :
    bitdata[287:283] == 5'b01100 ? cell_81_14 :
    bitdata[287:283] == 5'b11100 ? cell_81_15 :
    bitdata[287:283] == 5'b00010 ? cell_81_16 :
    bitdata[287:283] == 5'b10010 ? cell_81_17 :
    bitdata[287:283] == 5'b01010 ? cell_81_18 :
    bitdata[287:283] == 5'b11010 ? cell_81_19 :
    bitdata[287:283] == 5'b00110 ? cell_81_20 :
    bitdata[287:283] == 5'b10110 ? cell_81_21 :
    bitdata[287:283] == 5'b01110 ? cell_81_22 :
    bitdata[287:283] == 5'b11110 ? cell_81_23 :
    bitdata[287:283] == 5'b00001 ? cell_81_24 : 1'bx);
assign sw_0_0_25_up2 =
   (bitdata[292:288] == 5'b00000 ? cell_63_8 :
    bitdata[292:288] == 5'b10000 ? cell_63_9 :
    bitdata[292:288] == 5'b01000 ? cell_81_10 :
    bitdata[292:288] == 5'b11000 ? cell_81_11 :
    bitdata[292:288] == 5'b00100 ? cell_81_12 :
    bitdata[292:288] == 5'b10100 ? cell_81_13 :
    bitdata[292:288] == 5'b01100 ? cell_81_14 :
    bitdata[292:288] == 5'b11100 ? cell_81_15 :
    bitdata[292:288] == 5'b00010 ? cell_81_16 :
    bitdata[292:288] == 5'b10010 ? cell_81_17 :
    bitdata[292:288] == 5'b01010 ? cell_81_18 :
    bitdata[292:288] == 5'b11010 ? cell_81_19 :
    bitdata[292:288] == 5'b00110 ? cell_81_20 :
    bitdata[292:288] == 5'b10110 ? cell_81_21 :
    bitdata[292:288] == 5'b01110 ? cell_81_22 :
    bitdata[292:288] == 5'b11110 ? cell_81_23 :
    bitdata[292:288] == 5'b00001 ? cell_81_24 : 1'bx);
assign sw_0_0_25_up3 =
   (bitdata[297:293] == 5'b00000 ? cell_63_8 :
    bitdata[297:293] == 5'b10000 ? cell_63_9 :
    bitdata[297:293] == 5'b01000 ? cell_81_10 :
    bitdata[297:293] == 5'b11000 ? cell_81_11 :
    bitdata[297:293] == 5'b00100 ? cell_81_12 :
    bitdata[297:293] == 5'b10100 ? cell_81_13 :
    bitdata[297:293] == 5'b01100 ? cell_81_14 :
    bitdata[297:293] == 5'b11100 ? cell_81_15 :
    bitdata[297:293] == 5'b00010 ? cell_81_16 :
    bitdata[297:293] == 5'b10010 ? cell_81_17 :
    bitdata[297:293] == 5'b01010 ? cell_81_18 :
    bitdata[297:293] == 5'b11010 ? cell_81_19 :
    bitdata[297:293] == 5'b00110 ? cell_81_20 :
    bitdata[297:293] == 5'b10110 ? cell_81_21 :
    bitdata[297:293] == 5'b01110 ? cell_81_22 :
    bitdata[297:293] == 5'b11110 ? cell_81_23 :
    bitdata[297:293] == 5'b00001 ? cell_81_24 : 1'bx);
assign sw_0_0_26_down0 =
   (bitdata[91:89] == 3'b101 ? sw_0_0_7_down0 :
    bitdata[91:89] == 3'b000 ? sw_0_0_24_up0 :
    bitdata[91:89] == 3'b100 ? sw_0_0_25_up0 :
    bitdata[91:89] == 3'b010 ? sw_0_0_25_up1 :
    bitdata[91:89] == 3'b110 ? sw_0_0_25_up2 :
    bitdata[91:89] == 3'b001 ? sw_0_0_25_up3 : 1'bx);
assign sw_0_0_26_down1 =
   (bitdata[94:92] == 3'b101 ? sw_0_0_7_down0 :
    bitdata[94:92] == 3'b000 ? sw_0_0_24_up0 :
    bitdata[94:92] == 3'b100 ? sw_0_0_25_up0 :
    bitdata[94:92] == 3'b010 ? sw_0_0_25_up1 :
    bitdata[94:92] == 3'b110 ? sw_0_0_25_up2 :
    bitdata[94:92] == 3'b001 ? sw_0_0_25_up3 : 1'bx);
assign sw_0_0_26_up0 = cell_6_0;
assign sw_0_0_2_down0 = sw_0_0_1_up0;
assign sw_0_0_2_up0 =
   (bitdata[8:8] == 1'b0 ? sw_0_0_6_up0 :
    bitdata[8:8] == 1'b1 ? sw_0_0_7_up0 : 1'bx);
assign sw_0_0_3_down0 =
   (bitdata[3:2] == 2'b01 ? sw_0_0_1_down0 :
    bitdata[3:2] == 2'b00 ? sw_0_0_4_up0 :
    bitdata[3:2] == 2'b10 ? sw_0_0_5_up0 : 1'bx);
assign sw_0_0_3_up0 =
   (bitdata[14:11] == 4'b0000 ? sw_0_0_8_up0 :
    bitdata[14:11] == 4'b1000 ? sw_0_0_8_up1 :
    bitdata[14:11] == 4'b0100 ? sw_0_0_8_up2 :
    bitdata[14:11] == 4'b1100 ? sw_0_0_9_up0 :
    bitdata[14:11] == 4'b0010 ? sw_0_0_9_up1 :
    bitdata[14:11] == 4'b1010 ? sw_0_0_9_up2 :
    bitdata[14:11] == 4'b0110 ? sw_0_0_9_up3 :
    bitdata[14:11] == 4'b1110 ? sw_0_0_10_up0 :
    bitdata[14:11] == 4'b0001 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_4_down0 =
   (bitdata[5:4] == 2'b01 ? sw_0_0_1_down0 :
    bitdata[5:4] == 2'b00 ? sw_0_0_3_up0 :
    bitdata[5:4] == 2'b10 ? sw_0_0_5_up0 : 1'bx);
assign sw_0_0_4_up0 =
   (bitdata[50:50] == 1'b0 ? sw_0_0_12_up0 :
    bitdata[50:50] == 1'b1 ? sw_0_0_15_up0 : 1'bx);
assign sw_0_0_5_down0 =
   (bitdata[7:6] == 2'b01 ? sw_0_0_1_down0 :
    bitdata[7:6] == 2'b00 ? sw_0_0_3_up0 :
    bitdata[7:6] == 2'b10 ? sw_0_0_4_up0 : 1'bx);
assign sw_0_0_5_up0 =
   (bitdata[56:56] == 1'b0 ? sw_0_0_16_up0 :
    bitdata[56:56] == 1'b1 ? sw_0_0_18_up0 : 1'bx);
assign sw_0_0_6_down0 =
   (bitdata[9:9] == 1'b1 ? sw_0_0_2_down0 :
    bitdata[9:9] == 1'b0 ? sw_0_0_7_up0 : 1'bx);
assign sw_0_0_6_up0 =
   (bitdata[64:63] == 2'b00 ? sw_0_0_20_up0 :
    bitdata[64:63] == 2'b10 ? sw_0_0_22_up0 :
    bitdata[64:63] == 2'b01 ? sw_0_0_23_up0 : 1'bx);
assign sw_0_0_7_down0 =
   (bitdata[10:10] == 1'b1 ? sw_0_0_2_down0 :
    bitdata[10:10] == 1'b0 ? sw_0_0_6_up0 : 1'bx);
assign sw_0_0_7_up0 =
   (bitdata[73:71] == 3'b000 ? sw_0_0_24_up0 :
    bitdata[73:71] == 3'b100 ? sw_0_0_25_up0 :
    bitdata[73:71] == 3'b010 ? sw_0_0_25_up1 :
    bitdata[73:71] == 3'b110 ? sw_0_0_25_up2 :
    bitdata[73:71] == 3'b001 ? sw_0_0_25_up3 :
    bitdata[73:71] == 3'b101 ? sw_0_0_26_up0 : 1'bx);
assign sw_0_0_8_down0 =
   (bitdata[17:15] == 3'b011 ? sw_0_0_3_down0 :
    bitdata[17:15] == 3'b000 ? sw_0_0_9_up0 :
    bitdata[17:15] == 3'b100 ? sw_0_0_9_up1 :
    bitdata[17:15] == 3'b010 ? sw_0_0_9_up2 :
    bitdata[17:15] == 3'b110 ? sw_0_0_9_up3 :
    bitdata[17:15] == 3'b001 ? sw_0_0_10_up0 :
    bitdata[17:15] == 3'b101 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_8_down1 =
   (bitdata[20:18] == 3'b011 ? sw_0_0_3_down0 :
    bitdata[20:18] == 3'b000 ? sw_0_0_9_up0 :
    bitdata[20:18] == 3'b100 ? sw_0_0_9_up1 :
    bitdata[20:18] == 3'b010 ? sw_0_0_9_up2 :
    bitdata[20:18] == 3'b110 ? sw_0_0_9_up3 :
    bitdata[20:18] == 3'b001 ? sw_0_0_10_up0 :
    bitdata[20:18] == 3'b101 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_8_down2 =
   (bitdata[23:21] == 3'b011 ? sw_0_0_3_down0 :
    bitdata[23:21] == 3'b000 ? sw_0_0_9_up0 :
    bitdata[23:21] == 3'b100 ? sw_0_0_9_up1 :
    bitdata[23:21] == 3'b010 ? sw_0_0_9_up2 :
    bitdata[23:21] == 3'b110 ? sw_0_0_9_up3 :
    bitdata[23:21] == 3'b001 ? sw_0_0_10_up0 :
    bitdata[23:21] == 3'b101 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_8_down3 =
   (bitdata[26:24] == 3'b011 ? sw_0_0_3_down0 :
    bitdata[26:24] == 3'b000 ? sw_0_0_9_up0 :
    bitdata[26:24] == 3'b100 ? sw_0_0_9_up1 :
    bitdata[26:24] == 3'b010 ? sw_0_0_9_up2 :
    bitdata[26:24] == 3'b110 ? sw_0_0_9_up3 :
    bitdata[26:24] == 3'b001 ? sw_0_0_10_up0 :
    bitdata[26:24] == 3'b101 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_8_down4 =
   (bitdata[29:27] == 3'b011 ? sw_0_0_3_down0 :
    bitdata[29:27] == 3'b000 ? sw_0_0_9_up0 :
    bitdata[29:27] == 3'b100 ? sw_0_0_9_up1 :
    bitdata[29:27] == 3'b010 ? sw_0_0_9_up2 :
    bitdata[29:27] == 3'b110 ? sw_0_0_9_up3 :
    bitdata[29:27] == 3'b001 ? sw_0_0_10_up0 :
    bitdata[29:27] == 3'b101 ? sw_0_0_11_up0 : 1'bx);
assign sw_0_0_8_up0 =
   (bitdata[98:95] == 4'b0000 ? cell_61_6 :
    bitdata[98:95] == 4'b1000 ? cell_61_7 :
    bitdata[98:95] == 4'b0100 ? cell_71_5 :
    bitdata[98:95] == 4'b1100 ? cell_71_6 :
    bitdata[98:95] == 4'b0010 ? cell_71_7 :
    bitdata[98:95] == 4'b1010 ? cell_71_8 :
    bitdata[98:95] == 4'b0110 ? cell_80_6 :
    bitdata[98:95] == 4'b1110 ? cell_80_7 :
    bitdata[98:95] == 4'b0001 ? cell_80_8 :
    bitdata[98:95] == 4'b1001 ? cell_80_9 :
    bitdata[98:95] == 4'b0101 ? cell_80_10 :
    bitdata[98:95] == 4'b1101 ? cell_80_11 :
    bitdata[98:95] == 4'b0011 ? cell_80_12 :
    bitdata[98:95] == 4'b1011 ? cell_80_13 :
    bitdata[98:95] == 4'b0111 ? cell_80_14 :
    bitdata[98:95] == 4'b1111 ? cell_80_15 : 1'bx);
assign sw_0_0_8_up1 =
   (bitdata[102:99] == 4'b0000 ? cell_61_6 :
    bitdata[102:99] == 4'b1000 ? cell_61_7 :
    bitdata[102:99] == 4'b0100 ? cell_71_5 :
    bitdata[102:99] == 4'b1100 ? cell_71_6 :
    bitdata[102:99] == 4'b0010 ? cell_71_7 :
    bitdata[102:99] == 4'b1010 ? cell_71_8 :
    bitdata[102:99] == 4'b0110 ? cell_80_6 :
    bitdata[102:99] == 4'b1110 ? cell_80_7 :
    bitdata[102:99] == 4'b0001 ? cell_80_8 :
    bitdata[102:99] == 4'b1001 ? cell_80_9 :
    bitdata[102:99] == 4'b0101 ? cell_80_10 :
    bitdata[102:99] == 4'b1101 ? cell_80_11 :
    bitdata[102:99] == 4'b0011 ? cell_80_12 :
    bitdata[102:99] == 4'b1011 ? cell_80_13 :
    bitdata[102:99] == 4'b0111 ? cell_80_14 :
    bitdata[102:99] == 4'b1111 ? cell_80_15 : 1'bx);
assign sw_0_0_8_up2 =
   (bitdata[106:103] == 4'b0000 ? cell_61_6 :
    bitdata[106:103] == 4'b1000 ? cell_61_7 :
    bitdata[106:103] == 4'b0100 ? cell_71_5 :
    bitdata[106:103] == 4'b1100 ? cell_71_6 :
    bitdata[106:103] == 4'b0010 ? cell_71_7 :
    bitdata[106:103] == 4'b1010 ? cell_71_8 :
    bitdata[106:103] == 4'b0110 ? cell_80_6 :
    bitdata[106:103] == 4'b1110 ? cell_80_7 :
    bitdata[106:103] == 4'b0001 ? cell_80_8 :
    bitdata[106:103] == 4'b1001 ? cell_80_9 :
    bitdata[106:103] == 4'b0101 ? cell_80_10 :
    bitdata[106:103] == 4'b1101 ? cell_80_11 :
    bitdata[106:103] == 4'b0011 ? cell_80_12 :
    bitdata[106:103] == 4'b1011 ? cell_80_13 :
    bitdata[106:103] == 4'b0111 ? cell_80_14 :
    bitdata[106:103] == 4'b1111 ? cell_80_15 : 1'bx);
assign sw_0_0_9_up0 =
   (bitdata[167:166] == 2'b00 ? cell_0_0 :
    bitdata[167:166] == 2'b10 ? cell_14_0 :
    bitdata[167:166] == 2'b01 ? cell_45_0 :
    bitdata[167:166] == 2'b11 ? cell_82_0 : 1'bx);
assign sw_0_0_9_up1 =
   (bitdata[169:168] == 2'b00 ? cell_0_0 :
    bitdata[169:168] == 2'b10 ? cell_14_0 :
    bitdata[169:168] == 2'b01 ? cell_45_0 :
    bitdata[169:168] == 2'b11 ? cell_82_0 : 1'bx);
assign sw_0_0_9_up2 =
   (bitdata[171:170] == 2'b00 ? cell_0_0 :
    bitdata[171:170] == 2'b10 ? cell_14_0 :
    bitdata[171:170] == 2'b01 ? cell_45_0 :
    bitdata[171:170] == 2'b11 ? cell_82_0 : 1'bx);
assign sw_0_0_9_up3 =
   (bitdata[173:172] == 2'b00 ? cell_0_0 :
    bitdata[173:172] == 2'b10 ? cell_14_0 :
    bitdata[173:172] == 2'b01 ? cell_45_0 :
    bitdata[173:172] == 2'b11 ? cell_82_0 : 1'bx);
assign sw_0_1_10_down0 =
   (bitdata[479:475] == 5'b11110 ? sw_0_1_3_down0 :
    bitdata[479:475] == 5'b00001 ? sw_0_1_3_down1 :
    bitdata[479:475] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[479:475] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[479:475] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[479:475] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[479:475] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[479:475] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[479:475] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[479:475] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[479:475] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[479:475] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[479:475] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[479:475] == 5'b11010 ? sw_0_1_11_up0 :
    bitdata[479:475] == 5'b00110 ? sw_0_1_11_up1 :
    bitdata[479:475] == 5'b10110 ? sw_0_1_11_up2 :
    bitdata[479:475] == 5'b01110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_10_down1 =
   (bitdata[484:480] == 5'b11110 ? sw_0_1_3_down0 :
    bitdata[484:480] == 5'b00001 ? sw_0_1_3_down1 :
    bitdata[484:480] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[484:480] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[484:480] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[484:480] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[484:480] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[484:480] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[484:480] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[484:480] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[484:480] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[484:480] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[484:480] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[484:480] == 5'b11010 ? sw_0_1_11_up0 :
    bitdata[484:480] == 5'b00110 ? sw_0_1_11_up1 :
    bitdata[484:480] == 5'b10110 ? sw_0_1_11_up2 :
    bitdata[484:480] == 5'b01110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_10_down2 =
   (bitdata[489:485] == 5'b11110 ? sw_0_1_3_down0 :
    bitdata[489:485] == 5'b00001 ? sw_0_1_3_down1 :
    bitdata[489:485] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[489:485] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[489:485] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[489:485] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[489:485] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[489:485] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[489:485] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[489:485] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[489:485] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[489:485] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[489:485] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[489:485] == 5'b11010 ? sw_0_1_11_up0 :
    bitdata[489:485] == 5'b00110 ? sw_0_1_11_up1 :
    bitdata[489:485] == 5'b10110 ? sw_0_1_11_up2 :
    bitdata[489:485] == 5'b01110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_10_down3 =
   (bitdata[494:490] == 5'b11110 ? sw_0_1_3_down0 :
    bitdata[494:490] == 5'b00001 ? sw_0_1_3_down1 :
    bitdata[494:490] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[494:490] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[494:490] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[494:490] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[494:490] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[494:490] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[494:490] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[494:490] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[494:490] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[494:490] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[494:490] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[494:490] == 5'b11010 ? sw_0_1_11_up0 :
    bitdata[494:490] == 5'b00110 ? sw_0_1_11_up1 :
    bitdata[494:490] == 5'b10110 ? sw_0_1_11_up2 :
    bitdata[494:490] == 5'b01110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_10_down4 =
   (bitdata[499:495] == 5'b11110 ? sw_0_1_3_down0 :
    bitdata[499:495] == 5'b00001 ? sw_0_1_3_down1 :
    bitdata[499:495] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[499:495] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[499:495] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[499:495] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[499:495] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[499:495] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[499:495] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[499:495] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[499:495] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[499:495] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[499:495] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[499:495] == 5'b11010 ? sw_0_1_11_up0 :
    bitdata[499:495] == 5'b00110 ? sw_0_1_11_up1 :
    bitdata[499:495] == 5'b10110 ? sw_0_1_11_up2 :
    bitdata[499:495] == 5'b01110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_10_up0 =
   (bitdata[727:725] == 3'b000 ? cell_62_6 :
    bitdata[727:725] == 3'b100 ? cell_62_7 :
    bitdata[727:725] == 3'b010 ? cell_64_8 :
    bitdata[727:725] == 3'b110 ? cell_64_9 :
    bitdata[727:725] == 3'b001 ? cell_82_0 : 1'bx);
assign sw_0_1_10_up1 =
   (bitdata[730:728] == 3'b000 ? cell_62_6 :
    bitdata[730:728] == 3'b100 ? cell_62_7 :
    bitdata[730:728] == 3'b010 ? cell_64_8 :
    bitdata[730:728] == 3'b110 ? cell_64_9 :
    bitdata[730:728] == 3'b001 ? cell_82_0 : 1'bx);
assign sw_0_1_10_up2 =
   (bitdata[733:731] == 3'b000 ? cell_62_6 :
    bitdata[733:731] == 3'b100 ? cell_62_7 :
    bitdata[733:731] == 3'b010 ? cell_64_8 :
    bitdata[733:731] == 3'b110 ? cell_64_9 :
    bitdata[733:731] == 3'b001 ? cell_82_0 : 1'bx);
assign sw_0_1_11_down0 =
   (bitdata[503:500] == 4'b0111 ? sw_0_1_3_down0 :
    bitdata[503:500] == 4'b1111 ? sw_0_1_3_down1 :
    bitdata[503:500] == 4'b0000 ? sw_0_1_8_up0 :
    bitdata[503:500] == 4'b1000 ? sw_0_1_8_up1 :
    bitdata[503:500] == 4'b0100 ? sw_0_1_8_up2 :
    bitdata[503:500] == 4'b1100 ? sw_0_1_8_up3 :
    bitdata[503:500] == 4'b0010 ? sw_0_1_8_up4 :
    bitdata[503:500] == 4'b1010 ? sw_0_1_8_up5 :
    bitdata[503:500] == 4'b0110 ? sw_0_1_8_up6 :
    bitdata[503:500] == 4'b1110 ? sw_0_1_8_up7 :
    bitdata[503:500] == 4'b0001 ? sw_0_1_8_up8 :
    bitdata[503:500] == 4'b1001 ? sw_0_1_8_up9 :
    bitdata[503:500] == 4'b0101 ? sw_0_1_9_up0 :
    bitdata[503:500] == 4'b1101 ? sw_0_1_10_up0 :
    bitdata[503:500] == 4'b0011 ? sw_0_1_10_up1 :
    bitdata[503:500] == 4'b1011 ? sw_0_1_10_up2 : 1'bx);
assign sw_0_1_11_down1 =
   (bitdata[507:504] == 4'b0111 ? sw_0_1_3_down0 :
    bitdata[507:504] == 4'b1111 ? sw_0_1_3_down1 :
    bitdata[507:504] == 4'b0000 ? sw_0_1_8_up0 :
    bitdata[507:504] == 4'b1000 ? sw_0_1_8_up1 :
    bitdata[507:504] == 4'b0100 ? sw_0_1_8_up2 :
    bitdata[507:504] == 4'b1100 ? sw_0_1_8_up3 :
    bitdata[507:504] == 4'b0010 ? sw_0_1_8_up4 :
    bitdata[507:504] == 4'b1010 ? sw_0_1_8_up5 :
    bitdata[507:504] == 4'b0110 ? sw_0_1_8_up6 :
    bitdata[507:504] == 4'b1110 ? sw_0_1_8_up7 :
    bitdata[507:504] == 4'b0001 ? sw_0_1_8_up8 :
    bitdata[507:504] == 4'b1001 ? sw_0_1_8_up9 :
    bitdata[507:504] == 4'b0101 ? sw_0_1_9_up0 :
    bitdata[507:504] == 4'b1101 ? sw_0_1_10_up0 :
    bitdata[507:504] == 4'b0011 ? sw_0_1_10_up1 :
    bitdata[507:504] == 4'b1011 ? sw_0_1_10_up2 : 1'bx);
assign sw_0_1_11_down2 =
   (bitdata[511:508] == 4'b0111 ? sw_0_1_3_down0 :
    bitdata[511:508] == 4'b1111 ? sw_0_1_3_down1 :
    bitdata[511:508] == 4'b0000 ? sw_0_1_8_up0 :
    bitdata[511:508] == 4'b1000 ? sw_0_1_8_up1 :
    bitdata[511:508] == 4'b0100 ? sw_0_1_8_up2 :
    bitdata[511:508] == 4'b1100 ? sw_0_1_8_up3 :
    bitdata[511:508] == 4'b0010 ? sw_0_1_8_up4 :
    bitdata[511:508] == 4'b1010 ? sw_0_1_8_up5 :
    bitdata[511:508] == 4'b0110 ? sw_0_1_8_up6 :
    bitdata[511:508] == 4'b1110 ? sw_0_1_8_up7 :
    bitdata[511:508] == 4'b0001 ? sw_0_1_8_up8 :
    bitdata[511:508] == 4'b1001 ? sw_0_1_8_up9 :
    bitdata[511:508] == 4'b0101 ? sw_0_1_9_up0 :
    bitdata[511:508] == 4'b1101 ? sw_0_1_10_up0 :
    bitdata[511:508] == 4'b0011 ? sw_0_1_10_up1 :
    bitdata[511:508] == 4'b1011 ? sw_0_1_10_up2 : 1'bx);
assign sw_0_1_11_down3 =
   (bitdata[515:512] == 4'b0111 ? sw_0_1_3_down0 :
    bitdata[515:512] == 4'b1111 ? sw_0_1_3_down1 :
    bitdata[515:512] == 4'b0000 ? sw_0_1_8_up0 :
    bitdata[515:512] == 4'b1000 ? sw_0_1_8_up1 :
    bitdata[515:512] == 4'b0100 ? sw_0_1_8_up2 :
    bitdata[515:512] == 4'b1100 ? sw_0_1_8_up3 :
    bitdata[515:512] == 4'b0010 ? sw_0_1_8_up4 :
    bitdata[515:512] == 4'b1010 ? sw_0_1_8_up5 :
    bitdata[515:512] == 4'b0110 ? sw_0_1_8_up6 :
    bitdata[515:512] == 4'b1110 ? sw_0_1_8_up7 :
    bitdata[515:512] == 4'b0001 ? sw_0_1_8_up8 :
    bitdata[515:512] == 4'b1001 ? sw_0_1_8_up9 :
    bitdata[515:512] == 4'b0101 ? sw_0_1_9_up0 :
    bitdata[515:512] == 4'b1101 ? sw_0_1_10_up0 :
    bitdata[515:512] == 4'b0011 ? sw_0_1_10_up1 :
    bitdata[515:512] == 4'b1011 ? sw_0_1_10_up2 : 1'bx);
assign sw_0_1_11_up0 =
   (bitdata[773:770] == 4'b0000 ? cell_61_6 :
    bitdata[773:770] == 4'b1000 ? cell_61_7 :
    bitdata[773:770] == 4'b0100 ? cell_63_8 :
    bitdata[773:770] == 4'b1100 ? cell_63_9 :
    bitdata[773:770] == 4'b0010 ? cell_71_5 :
    bitdata[773:770] == 4'b1010 ? cell_71_6 :
    bitdata[773:770] == 4'b0110 ? cell_71_7 :
    bitdata[773:770] == 4'b1110 ? cell_71_8 :
    bitdata[773:770] == 4'b0001 ? cell_83_0 : 1'bx);
assign sw_0_1_11_up1 =
   (bitdata[777:774] == 4'b0000 ? cell_61_6 :
    bitdata[777:774] == 4'b1000 ? cell_61_7 :
    bitdata[777:774] == 4'b0100 ? cell_63_8 :
    bitdata[777:774] == 4'b1100 ? cell_63_9 :
    bitdata[777:774] == 4'b0010 ? cell_71_5 :
    bitdata[777:774] == 4'b1010 ? cell_71_6 :
    bitdata[777:774] == 4'b0110 ? cell_71_7 :
    bitdata[777:774] == 4'b1110 ? cell_71_8 :
    bitdata[777:774] == 4'b0001 ? cell_83_0 : 1'bx);
assign sw_0_1_11_up2 =
   (bitdata[781:778] == 4'b0000 ? cell_61_6 :
    bitdata[781:778] == 4'b1000 ? cell_61_7 :
    bitdata[781:778] == 4'b0100 ? cell_63_8 :
    bitdata[781:778] == 4'b1100 ? cell_63_9 :
    bitdata[781:778] == 4'b0010 ? cell_71_5 :
    bitdata[781:778] == 4'b1010 ? cell_71_6 :
    bitdata[781:778] == 4'b0110 ? cell_71_7 :
    bitdata[781:778] == 4'b1110 ? cell_71_8 :
    bitdata[781:778] == 4'b0001 ? cell_83_0 : 1'bx);
assign sw_0_1_11_up3 =
   (bitdata[785:782] == 4'b0000 ? cell_61_6 :
    bitdata[785:782] == 4'b1000 ? cell_61_7 :
    bitdata[785:782] == 4'b0100 ? cell_63_8 :
    bitdata[785:782] == 4'b1100 ? cell_63_9 :
    bitdata[785:782] == 4'b0010 ? cell_71_5 :
    bitdata[785:782] == 4'b1010 ? cell_71_6 :
    bitdata[785:782] == 4'b0110 ? cell_71_7 :
    bitdata[785:782] == 4'b1110 ? cell_71_8 :
    bitdata[785:782] == 4'b0001 ? cell_83_0 : 1'bx);
assign sw_0_1_12_down0 =
   (bitdata[517:516] == 2'b10 ? sw_0_1_4_down0 :
    bitdata[517:516] == 2'b01 ? sw_0_1_4_down1 :
    bitdata[517:516] == 2'b00 ? sw_0_1_15_up0 : 1'bx);
assign sw_0_1_12_down1 =
   (bitdata[519:518] == 2'b10 ? sw_0_1_4_down0 :
    bitdata[519:518] == 2'b01 ? sw_0_1_4_down1 :
    bitdata[519:518] == 2'b00 ? sw_0_1_15_up0 : 1'bx);
assign sw_0_1_13_down0 =
   (bitdata[521:520] == 2'b10 ? sw_0_1_4_down0 :
    bitdata[521:520] == 2'b01 ? sw_0_1_4_down1 :
    bitdata[521:520] == 2'b00 ? sw_0_1_15_up0 : 1'bx);
assign sw_0_1_14_down0 =
   (bitdata[523:522] == 2'b10 ? sw_0_1_4_down0 :
    bitdata[523:522] == 2'b01 ? sw_0_1_4_down1 :
    bitdata[523:522] == 2'b00 ? sw_0_1_15_up0 : 1'bx);
assign sw_0_1_15_up0 =
   (bitdata[847:846] == 2'b00 ? cell_49_0 :
    bitdata[847:846] == 2'b10 ? cell_50_0 :
    bitdata[847:846] == 2'b01 ? cell_51_0 :
    bitdata[847:846] == 2'b11 ? cell_52_0 : 1'bx);
assign sw_0_1_16_up0 =
   (bitdata[849:848] == 2'b00 ? cell_45_0 :
    bitdata[849:848] == 2'b10 ? cell_46_0 :
    bitdata[849:848] == 2'b01 ? cell_47_0 :
    bitdata[849:848] == 2'b11 ? cell_48_0 : 1'bx);
assign sw_0_1_16_up1 =
   (bitdata[851:850] == 2'b00 ? cell_45_0 :
    bitdata[851:850] == 2'b10 ? cell_46_0 :
    bitdata[851:850] == 2'b01 ? cell_47_0 :
    bitdata[851:850] == 2'b11 ? cell_48_0 : 1'bx);
assign sw_0_1_17_down0 =
   (bitdata[533:530] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[533:530] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[533:530] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[533:530] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[533:530] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[533:530] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[533:530] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[533:530] == 4'b0100 ? sw_0_1_18_up0 :
    bitdata[533:530] == 4'b1100 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_17_down1 =
   (bitdata[537:534] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[537:534] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[537:534] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[537:534] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[537:534] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[537:534] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[537:534] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[537:534] == 4'b0100 ? sw_0_1_18_up0 :
    bitdata[537:534] == 4'b1100 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_17_down2 =
   (bitdata[541:538] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[541:538] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[541:538] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[541:538] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[541:538] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[541:538] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[541:538] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[541:538] == 4'b0100 ? sw_0_1_18_up0 :
    bitdata[541:538] == 4'b1100 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_17_up0 = cell_39_0;
assign sw_0_1_18_down0 =
   (bitdata[545:542] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[545:542] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[545:542] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[545:542] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[545:542] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[545:542] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[545:542] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[545:542] == 4'b0100 ? sw_0_1_17_up0 :
    bitdata[545:542] == 4'b1100 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_18_down1 =
   (bitdata[549:546] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[549:546] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[549:546] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[549:546] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[549:546] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[549:546] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[549:546] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[549:546] == 4'b0100 ? sw_0_1_17_up0 :
    bitdata[549:546] == 4'b1100 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_18_down2 =
   (bitdata[553:550] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[553:550] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[553:550] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[553:550] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[553:550] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[553:550] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[553:550] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[553:550] == 4'b0100 ? sw_0_1_17_up0 :
    bitdata[553:550] == 4'b1100 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_18_up0 =
   (bitdata[862:861] == 2'b00 ? cell_72_5 :
    bitdata[862:861] == 2'b10 ? cell_72_6 :
    bitdata[862:861] == 2'b01 ? cell_72_7 :
    bitdata[862:861] == 2'b11 ? cell_72_8 : 1'bx);
assign sw_0_1_19_down0 =
   (bitdata[557:554] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[557:554] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[557:554] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[557:554] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[557:554] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[557:554] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[557:554] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[557:554] == 4'b0100 ? sw_0_1_17_up0 :
    bitdata[557:554] == 4'b1100 ? sw_0_1_18_up0 : 1'bx);
assign sw_0_1_19_down1 =
   (bitdata[561:558] == 4'b0010 ? sw_0_1_5_down0 :
    bitdata[561:558] == 4'b1010 ? sw_0_1_5_down1 :
    bitdata[561:558] == 4'b0110 ? sw_0_1_5_down2 :
    bitdata[561:558] == 4'b1110 ? sw_0_1_5_down3 :
    bitdata[561:558] == 4'b0001 ? sw_0_1_5_down4 :
    bitdata[561:558] == 4'b0000 ? sw_0_1_16_up0 :
    bitdata[561:558] == 4'b1000 ? sw_0_1_16_up1 :
    bitdata[561:558] == 4'b0100 ? sw_0_1_17_up0 :
    bitdata[561:558] == 4'b1100 ? sw_0_1_18_up0 : 1'bx);
assign sw_0_1_19_up0 = cell_40_0;
assign sw_0_1_1_down0 = sw_0_1_2_up0;
assign sw_0_1_1_up0 =
   (bitdata[375:372] == 4'b0000 ? sw_0_1_3_up0 :
    bitdata[375:372] == 4'b1000 ? sw_0_1_3_up1 :
    bitdata[375:372] == 4'b0100 ? sw_0_1_3_up2 :
    bitdata[375:372] == 4'b1100 ? sw_0_1_3_up3 :
    bitdata[375:372] == 4'b0010 ? sw_0_1_3_up4 :
    bitdata[375:372] == 4'b1010 ? sw_0_1_3_up5 :
    bitdata[375:372] == 4'b0110 ? sw_0_1_4_up0 :
    bitdata[375:372] == 4'b1110 ? sw_0_1_5_up0 :
    bitdata[375:372] == 4'b0001 ? sw_0_1_5_up1 : 1'bx);
assign sw_0_1_20_down0 =
   (bitdata[564:563] == 2'b01 ? sw_0_1_6_down0 :
    bitdata[564:563] == 2'b00 ? sw_0_1_22_up0 :
    bitdata[564:563] == 2'b10 ? sw_0_1_23_up0 : 1'bx);
assign sw_0_1_21_down0 =
   (bitdata[566:565] == 2'b01 ? sw_0_1_6_down0 :
    bitdata[566:565] == 2'b00 ? sw_0_1_22_up0 :
    bitdata[566:565] == 2'b10 ? sw_0_1_23_up0 : 1'bx);
assign sw_0_1_22_down0 =
   (bitdata[567:567] == 1'b1 ? sw_0_1_6_down0 :
    bitdata[567:567] == 1'b0 ? sw_0_1_23_up0 : 1'bx);
assign sw_0_1_22_up0 =
   (bitdata[891:890] == 2'b00 ? cell_19_0 :
    bitdata[891:890] == 2'b10 ? cell_20_0 :
    bitdata[891:890] == 2'b01 ? cell_21_0 : 1'bx);
assign sw_0_1_23_up0 =
   (bitdata[896:895] == 2'b00 ? cell_15_0 :
    bitdata[896:895] == 2'b10 ? cell_16_0 :
    bitdata[896:895] == 2'b01 ? cell_17_0 :
    bitdata[896:895] == 2'b11 ? cell_18_0 : 1'bx);
assign sw_0_1_24_down0 =
   (bitdata[571:570] == 2'b01 ? sw_0_1_7_down0 :
    bitdata[571:570] == 2'b00 ? sw_0_1_25_up0 :
    bitdata[571:570] == 2'b10 ? sw_0_1_26_up0 : 1'bx);
assign sw_0_1_24_up0 = cell_14_0;
assign sw_0_1_25_down0 =
   (bitdata[573:572] == 2'b01 ? sw_0_1_7_down0 :
    bitdata[573:572] == 2'b00 ? sw_0_1_24_up0 :
    bitdata[573:572] == 2'b10 ? sw_0_1_26_up0 : 1'bx);
assign sw_0_1_25_up0 =
   (bitdata[904:903] == 2'b00 ? cell_6_0 :
    bitdata[904:903] == 2'b10 ? cell_7_0 :
    bitdata[904:903] == 2'b01 ? cell_8_0 : 1'bx);
assign sw_0_1_26_down0 =
   (bitdata[575:574] == 2'b01 ? sw_0_1_7_down0 :
    bitdata[575:574] == 2'b00 ? sw_0_1_24_up0 :
    bitdata[575:574] == 2'b10 ? sw_0_1_25_up0 : 1'bx);
assign sw_0_1_26_up0 =
   (bitdata[908:908] == 1'b0 ? cell_0_0 :
    bitdata[908:908] == 1'b1 ? cell_3_0 : 1'bx);
assign sw_0_1_2_down0 = sw_0_1_1_up0;
assign sw_0_1_2_up0 =
   (bitdata[403:403] == 1'b0 ? sw_0_1_6_up0 :
    bitdata[403:403] == 1'b1 ? sw_0_1_7_up0 : 1'bx);
assign sw_0_1_3_down0 =
   (bitdata[377:376] == 2'b11 ? sw_0_1_1_down0 :
    bitdata[377:376] == 2'b00 ? sw_0_1_4_up0 :
    bitdata[377:376] == 2'b10 ? sw_0_1_5_up0 :
    bitdata[377:376] == 2'b01 ? sw_0_1_5_up1 : 1'bx);
assign sw_0_1_3_down1 =
   (bitdata[379:378] == 2'b11 ? sw_0_1_1_down0 :
    bitdata[379:378] == 2'b00 ? sw_0_1_4_up0 :
    bitdata[379:378] == 2'b10 ? sw_0_1_5_up0 :
    bitdata[379:378] == 2'b01 ? sw_0_1_5_up1 : 1'bx);
assign sw_0_1_3_up0 =
   (bitdata[410:406] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[410:406] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[410:406] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[410:406] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[410:406] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[410:406] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[410:406] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[410:406] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[410:406] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[410:406] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[410:406] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[410:406] == 5'b11010 ? sw_0_1_10_up0 :
    bitdata[410:406] == 5'b00110 ? sw_0_1_10_up1 :
    bitdata[410:406] == 5'b10110 ? sw_0_1_10_up2 :
    bitdata[410:406] == 5'b01110 ? sw_0_1_11_up0 :
    bitdata[410:406] == 5'b11110 ? sw_0_1_11_up1 :
    bitdata[410:406] == 5'b00001 ? sw_0_1_11_up2 :
    bitdata[410:406] == 5'b10001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_3_up1 =
   (bitdata[415:411] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[415:411] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[415:411] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[415:411] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[415:411] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[415:411] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[415:411] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[415:411] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[415:411] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[415:411] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[415:411] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[415:411] == 5'b11010 ? sw_0_1_10_up0 :
    bitdata[415:411] == 5'b00110 ? sw_0_1_10_up1 :
    bitdata[415:411] == 5'b10110 ? sw_0_1_10_up2 :
    bitdata[415:411] == 5'b01110 ? sw_0_1_11_up0 :
    bitdata[415:411] == 5'b11110 ? sw_0_1_11_up1 :
    bitdata[415:411] == 5'b00001 ? sw_0_1_11_up2 :
    bitdata[415:411] == 5'b10001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_3_up2 =
   (bitdata[420:416] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[420:416] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[420:416] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[420:416] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[420:416] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[420:416] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[420:416] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[420:416] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[420:416] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[420:416] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[420:416] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[420:416] == 5'b11010 ? sw_0_1_10_up0 :
    bitdata[420:416] == 5'b00110 ? sw_0_1_10_up1 :
    bitdata[420:416] == 5'b10110 ? sw_0_1_10_up2 :
    bitdata[420:416] == 5'b01110 ? sw_0_1_11_up0 :
    bitdata[420:416] == 5'b11110 ? sw_0_1_11_up1 :
    bitdata[420:416] == 5'b00001 ? sw_0_1_11_up2 :
    bitdata[420:416] == 5'b10001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_3_up3 =
   (bitdata[425:421] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[425:421] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[425:421] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[425:421] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[425:421] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[425:421] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[425:421] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[425:421] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[425:421] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[425:421] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[425:421] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[425:421] == 5'b11010 ? sw_0_1_10_up0 :
    bitdata[425:421] == 5'b00110 ? sw_0_1_10_up1 :
    bitdata[425:421] == 5'b10110 ? sw_0_1_10_up2 :
    bitdata[425:421] == 5'b01110 ? sw_0_1_11_up0 :
    bitdata[425:421] == 5'b11110 ? sw_0_1_11_up1 :
    bitdata[425:421] == 5'b00001 ? sw_0_1_11_up2 :
    bitdata[425:421] == 5'b10001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_3_up4 =
   (bitdata[430:426] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[430:426] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[430:426] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[430:426] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[430:426] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[430:426] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[430:426] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[430:426] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[430:426] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[430:426] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[430:426] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[430:426] == 5'b11010 ? sw_0_1_10_up0 :
    bitdata[430:426] == 5'b00110 ? sw_0_1_10_up1 :
    bitdata[430:426] == 5'b10110 ? sw_0_1_10_up2 :
    bitdata[430:426] == 5'b01110 ? sw_0_1_11_up0 :
    bitdata[430:426] == 5'b11110 ? sw_0_1_11_up1 :
    bitdata[430:426] == 5'b00001 ? sw_0_1_11_up2 :
    bitdata[430:426] == 5'b10001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_3_up5 =
   (bitdata[435:431] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[435:431] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[435:431] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[435:431] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[435:431] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[435:431] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[435:431] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[435:431] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[435:431] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[435:431] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[435:431] == 5'b01010 ? sw_0_1_9_up0 :
    bitdata[435:431] == 5'b11010 ? sw_0_1_10_up0 :
    bitdata[435:431] == 5'b00110 ? sw_0_1_10_up1 :
    bitdata[435:431] == 5'b10110 ? sw_0_1_10_up2 :
    bitdata[435:431] == 5'b01110 ? sw_0_1_11_up0 :
    bitdata[435:431] == 5'b11110 ? sw_0_1_11_up1 :
    bitdata[435:431] == 5'b00001 ? sw_0_1_11_up2 :
    bitdata[435:431] == 5'b10001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_4_down0 =
   (bitdata[383:380] == 4'b0001 ? sw_0_1_1_down0 :
    bitdata[383:380] == 4'b0000 ? sw_0_1_3_up0 :
    bitdata[383:380] == 4'b1000 ? sw_0_1_3_up1 :
    bitdata[383:380] == 4'b0100 ? sw_0_1_3_up2 :
    bitdata[383:380] == 4'b1100 ? sw_0_1_3_up3 :
    bitdata[383:380] == 4'b0010 ? sw_0_1_3_up4 :
    bitdata[383:380] == 4'b1010 ? sw_0_1_3_up5 :
    bitdata[383:380] == 4'b0110 ? sw_0_1_5_up0 :
    bitdata[383:380] == 4'b1110 ? sw_0_1_5_up1 : 1'bx);
assign sw_0_1_4_down1 =
   (bitdata[387:384] == 4'b0001 ? sw_0_1_1_down0 :
    bitdata[387:384] == 4'b0000 ? sw_0_1_3_up0 :
    bitdata[387:384] == 4'b1000 ? sw_0_1_3_up1 :
    bitdata[387:384] == 4'b0100 ? sw_0_1_3_up2 :
    bitdata[387:384] == 4'b1100 ? sw_0_1_3_up3 :
    bitdata[387:384] == 4'b0010 ? sw_0_1_3_up4 :
    bitdata[387:384] == 4'b1010 ? sw_0_1_3_up5 :
    bitdata[387:384] == 4'b0110 ? sw_0_1_5_up0 :
    bitdata[387:384] == 4'b1110 ? sw_0_1_5_up1 : 1'bx);
assign sw_0_1_4_up0 = sw_0_1_15_up0;
assign sw_0_1_5_down0 =
   (bitdata[390:388] == 3'b111 ? sw_0_1_1_down0 :
    bitdata[390:388] == 3'b000 ? sw_0_1_3_up0 :
    bitdata[390:388] == 3'b100 ? sw_0_1_3_up1 :
    bitdata[390:388] == 3'b010 ? sw_0_1_3_up2 :
    bitdata[390:388] == 3'b110 ? sw_0_1_3_up3 :
    bitdata[390:388] == 3'b001 ? sw_0_1_3_up4 :
    bitdata[390:388] == 3'b101 ? sw_0_1_3_up5 :
    bitdata[390:388] == 3'b011 ? sw_0_1_4_up0 : 1'bx);
assign sw_0_1_5_down1 =
   (bitdata[393:391] == 3'b111 ? sw_0_1_1_down0 :
    bitdata[393:391] == 3'b000 ? sw_0_1_3_up0 :
    bitdata[393:391] == 3'b100 ? sw_0_1_3_up1 :
    bitdata[393:391] == 3'b010 ? sw_0_1_3_up2 :
    bitdata[393:391] == 3'b110 ? sw_0_1_3_up3 :
    bitdata[393:391] == 3'b001 ? sw_0_1_3_up4 :
    bitdata[393:391] == 3'b101 ? sw_0_1_3_up5 :
    bitdata[393:391] == 3'b011 ? sw_0_1_4_up0 : 1'bx);
assign sw_0_1_5_down2 =
   (bitdata[396:394] == 3'b111 ? sw_0_1_1_down0 :
    bitdata[396:394] == 3'b000 ? sw_0_1_3_up0 :
    bitdata[396:394] == 3'b100 ? sw_0_1_3_up1 :
    bitdata[396:394] == 3'b010 ? sw_0_1_3_up2 :
    bitdata[396:394] == 3'b110 ? sw_0_1_3_up3 :
    bitdata[396:394] == 3'b001 ? sw_0_1_3_up4 :
    bitdata[396:394] == 3'b101 ? sw_0_1_3_up5 :
    bitdata[396:394] == 3'b011 ? sw_0_1_4_up0 : 1'bx);
assign sw_0_1_5_down3 =
   (bitdata[399:397] == 3'b111 ? sw_0_1_1_down0 :
    bitdata[399:397] == 3'b000 ? sw_0_1_3_up0 :
    bitdata[399:397] == 3'b100 ? sw_0_1_3_up1 :
    bitdata[399:397] == 3'b010 ? sw_0_1_3_up2 :
    bitdata[399:397] == 3'b110 ? sw_0_1_3_up3 :
    bitdata[399:397] == 3'b001 ? sw_0_1_3_up4 :
    bitdata[399:397] == 3'b101 ? sw_0_1_3_up5 :
    bitdata[399:397] == 3'b011 ? sw_0_1_4_up0 : 1'bx);
assign sw_0_1_5_down4 =
   (bitdata[402:400] == 3'b111 ? sw_0_1_1_down0 :
    bitdata[402:400] == 3'b000 ? sw_0_1_3_up0 :
    bitdata[402:400] == 3'b100 ? sw_0_1_3_up1 :
    bitdata[402:400] == 3'b010 ? sw_0_1_3_up2 :
    bitdata[402:400] == 3'b110 ? sw_0_1_3_up3 :
    bitdata[402:400] == 3'b001 ? sw_0_1_3_up4 :
    bitdata[402:400] == 3'b101 ? sw_0_1_3_up5 :
    bitdata[402:400] == 3'b011 ? sw_0_1_4_up0 : 1'bx);
assign sw_0_1_5_up0 =
   (bitdata[526:524] == 3'b000 ? sw_0_1_16_up0 :
    bitdata[526:524] == 3'b100 ? sw_0_1_16_up1 :
    bitdata[526:524] == 3'b010 ? sw_0_1_17_up0 :
    bitdata[526:524] == 3'b110 ? sw_0_1_18_up0 :
    bitdata[526:524] == 3'b001 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_5_up1 =
   (bitdata[529:527] == 3'b000 ? sw_0_1_16_up0 :
    bitdata[529:527] == 3'b100 ? sw_0_1_16_up1 :
    bitdata[529:527] == 3'b010 ? sw_0_1_17_up0 :
    bitdata[529:527] == 3'b110 ? sw_0_1_18_up0 :
    bitdata[529:527] == 3'b001 ? sw_0_1_19_up0 : 1'bx);
assign sw_0_1_6_down0 =
   (bitdata[404:404] == 1'b1 ? sw_0_1_2_down0 :
    bitdata[404:404] == 1'b0 ? sw_0_1_7_up0 : 1'bx);
assign sw_0_1_6_up0 =
   (bitdata[562:562] == 1'b0 ? sw_0_1_22_up0 :
    bitdata[562:562] == 1'b1 ? sw_0_1_23_up0 : 1'bx);
assign sw_0_1_7_down0 =
   (bitdata[405:405] == 1'b1 ? sw_0_1_2_down0 :
    bitdata[405:405] == 1'b0 ? sw_0_1_6_up0 : 1'bx);
assign sw_0_1_7_up0 =
   (bitdata[569:568] == 2'b00 ? sw_0_1_24_up0 :
    bitdata[569:568] == 2'b10 ? sw_0_1_25_up0 :
    bitdata[569:568] == 2'b01 ? sw_0_1_26_up0 : 1'bx);
assign sw_0_1_8_down0 =
   (bitdata[439:436] == 4'b0001 ? sw_0_1_3_down0 :
    bitdata[439:436] == 4'b1001 ? sw_0_1_3_down1 :
    bitdata[439:436] == 4'b0000 ? sw_0_1_9_up0 :
    bitdata[439:436] == 4'b1000 ? sw_0_1_10_up0 :
    bitdata[439:436] == 4'b0100 ? sw_0_1_10_up1 :
    bitdata[439:436] == 4'b1100 ? sw_0_1_10_up2 :
    bitdata[439:436] == 4'b0010 ? sw_0_1_11_up0 :
    bitdata[439:436] == 4'b1010 ? sw_0_1_11_up1 :
    bitdata[439:436] == 4'b0110 ? sw_0_1_11_up2 :
    bitdata[439:436] == 4'b1110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_8_down1 =
   (bitdata[443:440] == 4'b0001 ? sw_0_1_3_down0 :
    bitdata[443:440] == 4'b1001 ? sw_0_1_3_down1 :
    bitdata[443:440] == 4'b0000 ? sw_0_1_9_up0 :
    bitdata[443:440] == 4'b1000 ? sw_0_1_10_up0 :
    bitdata[443:440] == 4'b0100 ? sw_0_1_10_up1 :
    bitdata[443:440] == 4'b1100 ? sw_0_1_10_up2 :
    bitdata[443:440] == 4'b0010 ? sw_0_1_11_up0 :
    bitdata[443:440] == 4'b1010 ? sw_0_1_11_up1 :
    bitdata[443:440] == 4'b0110 ? sw_0_1_11_up2 :
    bitdata[443:440] == 4'b1110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_8_down2 =
   (bitdata[447:444] == 4'b0001 ? sw_0_1_3_down0 :
    bitdata[447:444] == 4'b1001 ? sw_0_1_3_down1 :
    bitdata[447:444] == 4'b0000 ? sw_0_1_9_up0 :
    bitdata[447:444] == 4'b1000 ? sw_0_1_10_up0 :
    bitdata[447:444] == 4'b0100 ? sw_0_1_10_up1 :
    bitdata[447:444] == 4'b1100 ? sw_0_1_10_up2 :
    bitdata[447:444] == 4'b0010 ? sw_0_1_11_up0 :
    bitdata[447:444] == 4'b1010 ? sw_0_1_11_up1 :
    bitdata[447:444] == 4'b0110 ? sw_0_1_11_up2 :
    bitdata[447:444] == 4'b1110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_8_down3 =
   (bitdata[451:448] == 4'b0001 ? sw_0_1_3_down0 :
    bitdata[451:448] == 4'b1001 ? sw_0_1_3_down1 :
    bitdata[451:448] == 4'b0000 ? sw_0_1_9_up0 :
    bitdata[451:448] == 4'b1000 ? sw_0_1_10_up0 :
    bitdata[451:448] == 4'b0100 ? sw_0_1_10_up1 :
    bitdata[451:448] == 4'b1100 ? sw_0_1_10_up2 :
    bitdata[451:448] == 4'b0010 ? sw_0_1_11_up0 :
    bitdata[451:448] == 4'b1010 ? sw_0_1_11_up1 :
    bitdata[451:448] == 4'b0110 ? sw_0_1_11_up2 :
    bitdata[451:448] == 4'b1110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_8_down4 =
   (bitdata[455:452] == 4'b0001 ? sw_0_1_3_down0 :
    bitdata[455:452] == 4'b1001 ? sw_0_1_3_down1 :
    bitdata[455:452] == 4'b0000 ? sw_0_1_9_up0 :
    bitdata[455:452] == 4'b1000 ? sw_0_1_10_up0 :
    bitdata[455:452] == 4'b0100 ? sw_0_1_10_up1 :
    bitdata[455:452] == 4'b1100 ? sw_0_1_10_up2 :
    bitdata[455:452] == 4'b0010 ? sw_0_1_11_up0 :
    bitdata[455:452] == 4'b1010 ? sw_0_1_11_up1 :
    bitdata[455:452] == 4'b0110 ? sw_0_1_11_up2 :
    bitdata[455:452] == 4'b1110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_8_down5 =
   (bitdata[459:456] == 4'b0001 ? sw_0_1_3_down0 :
    bitdata[459:456] == 4'b1001 ? sw_0_1_3_down1 :
    bitdata[459:456] == 4'b0000 ? sw_0_1_9_up0 :
    bitdata[459:456] == 4'b1000 ? sw_0_1_10_up0 :
    bitdata[459:456] == 4'b0100 ? sw_0_1_10_up1 :
    bitdata[459:456] == 4'b1100 ? sw_0_1_10_up2 :
    bitdata[459:456] == 4'b0010 ? sw_0_1_11_up0 :
    bitdata[459:456] == 4'b1010 ? sw_0_1_11_up1 :
    bitdata[459:456] == 4'b0110 ? sw_0_1_11_up2 :
    bitdata[459:456] == 4'b1110 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_8_up0 =
   (bitdata[580:576] == 5'b00000 ? cell_80_6 :
    bitdata[580:576] == 5'b10000 ? cell_80_7 :
    bitdata[580:576] == 5'b01000 ? cell_80_8 :
    bitdata[580:576] == 5'b11000 ? cell_80_9 :
    bitdata[580:576] == 5'b00100 ? cell_80_10 :
    bitdata[580:576] == 5'b10100 ? cell_80_11 :
    bitdata[580:576] == 5'b01100 ? cell_80_12 :
    bitdata[580:576] == 5'b11100 ? cell_80_13 :
    bitdata[580:576] == 5'b00010 ? cell_80_14 :
    bitdata[580:576] == 5'b10010 ? cell_80_15 :
    bitdata[580:576] == 5'b01010 ? cell_81_10 :
    bitdata[580:576] == 5'b11010 ? cell_81_11 :
    bitdata[580:576] == 5'b00110 ? cell_81_12 :
    bitdata[580:576] == 5'b10110 ? cell_81_13 :
    bitdata[580:576] == 5'b01110 ? cell_81_14 :
    bitdata[580:576] == 5'b11110 ? cell_81_15 :
    bitdata[580:576] == 5'b00001 ? cell_81_16 :
    bitdata[580:576] == 5'b10001 ? cell_81_17 :
    bitdata[580:576] == 5'b01001 ? cell_81_18 :
    bitdata[580:576] == 5'b11001 ? cell_81_19 :
    bitdata[580:576] == 5'b00101 ? cell_81_20 :
    bitdata[580:576] == 5'b10101 ? cell_81_21 :
    bitdata[580:576] == 5'b01101 ? cell_81_22 :
    bitdata[580:576] == 5'b11101 ? cell_81_23 :
    bitdata[580:576] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up1 =
   (bitdata[585:581] == 5'b00000 ? cell_80_6 :
    bitdata[585:581] == 5'b10000 ? cell_80_7 :
    bitdata[585:581] == 5'b01000 ? cell_80_8 :
    bitdata[585:581] == 5'b11000 ? cell_80_9 :
    bitdata[585:581] == 5'b00100 ? cell_80_10 :
    bitdata[585:581] == 5'b10100 ? cell_80_11 :
    bitdata[585:581] == 5'b01100 ? cell_80_12 :
    bitdata[585:581] == 5'b11100 ? cell_80_13 :
    bitdata[585:581] == 5'b00010 ? cell_80_14 :
    bitdata[585:581] == 5'b10010 ? cell_80_15 :
    bitdata[585:581] == 5'b01010 ? cell_81_10 :
    bitdata[585:581] == 5'b11010 ? cell_81_11 :
    bitdata[585:581] == 5'b00110 ? cell_81_12 :
    bitdata[585:581] == 5'b10110 ? cell_81_13 :
    bitdata[585:581] == 5'b01110 ? cell_81_14 :
    bitdata[585:581] == 5'b11110 ? cell_81_15 :
    bitdata[585:581] == 5'b00001 ? cell_81_16 :
    bitdata[585:581] == 5'b10001 ? cell_81_17 :
    bitdata[585:581] == 5'b01001 ? cell_81_18 :
    bitdata[585:581] == 5'b11001 ? cell_81_19 :
    bitdata[585:581] == 5'b00101 ? cell_81_20 :
    bitdata[585:581] == 5'b10101 ? cell_81_21 :
    bitdata[585:581] == 5'b01101 ? cell_81_22 :
    bitdata[585:581] == 5'b11101 ? cell_81_23 :
    bitdata[585:581] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up2 =
   (bitdata[590:586] == 5'b00000 ? cell_80_6 :
    bitdata[590:586] == 5'b10000 ? cell_80_7 :
    bitdata[590:586] == 5'b01000 ? cell_80_8 :
    bitdata[590:586] == 5'b11000 ? cell_80_9 :
    bitdata[590:586] == 5'b00100 ? cell_80_10 :
    bitdata[590:586] == 5'b10100 ? cell_80_11 :
    bitdata[590:586] == 5'b01100 ? cell_80_12 :
    bitdata[590:586] == 5'b11100 ? cell_80_13 :
    bitdata[590:586] == 5'b00010 ? cell_80_14 :
    bitdata[590:586] == 5'b10010 ? cell_80_15 :
    bitdata[590:586] == 5'b01010 ? cell_81_10 :
    bitdata[590:586] == 5'b11010 ? cell_81_11 :
    bitdata[590:586] == 5'b00110 ? cell_81_12 :
    bitdata[590:586] == 5'b10110 ? cell_81_13 :
    bitdata[590:586] == 5'b01110 ? cell_81_14 :
    bitdata[590:586] == 5'b11110 ? cell_81_15 :
    bitdata[590:586] == 5'b00001 ? cell_81_16 :
    bitdata[590:586] == 5'b10001 ? cell_81_17 :
    bitdata[590:586] == 5'b01001 ? cell_81_18 :
    bitdata[590:586] == 5'b11001 ? cell_81_19 :
    bitdata[590:586] == 5'b00101 ? cell_81_20 :
    bitdata[590:586] == 5'b10101 ? cell_81_21 :
    bitdata[590:586] == 5'b01101 ? cell_81_22 :
    bitdata[590:586] == 5'b11101 ? cell_81_23 :
    bitdata[590:586] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up3 =
   (bitdata[595:591] == 5'b00000 ? cell_80_6 :
    bitdata[595:591] == 5'b10000 ? cell_80_7 :
    bitdata[595:591] == 5'b01000 ? cell_80_8 :
    bitdata[595:591] == 5'b11000 ? cell_80_9 :
    bitdata[595:591] == 5'b00100 ? cell_80_10 :
    bitdata[595:591] == 5'b10100 ? cell_80_11 :
    bitdata[595:591] == 5'b01100 ? cell_80_12 :
    bitdata[595:591] == 5'b11100 ? cell_80_13 :
    bitdata[595:591] == 5'b00010 ? cell_80_14 :
    bitdata[595:591] == 5'b10010 ? cell_80_15 :
    bitdata[595:591] == 5'b01010 ? cell_81_10 :
    bitdata[595:591] == 5'b11010 ? cell_81_11 :
    bitdata[595:591] == 5'b00110 ? cell_81_12 :
    bitdata[595:591] == 5'b10110 ? cell_81_13 :
    bitdata[595:591] == 5'b01110 ? cell_81_14 :
    bitdata[595:591] == 5'b11110 ? cell_81_15 :
    bitdata[595:591] == 5'b00001 ? cell_81_16 :
    bitdata[595:591] == 5'b10001 ? cell_81_17 :
    bitdata[595:591] == 5'b01001 ? cell_81_18 :
    bitdata[595:591] == 5'b11001 ? cell_81_19 :
    bitdata[595:591] == 5'b00101 ? cell_81_20 :
    bitdata[595:591] == 5'b10101 ? cell_81_21 :
    bitdata[595:591] == 5'b01101 ? cell_81_22 :
    bitdata[595:591] == 5'b11101 ? cell_81_23 :
    bitdata[595:591] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up4 =
   (bitdata[600:596] == 5'b00000 ? cell_80_6 :
    bitdata[600:596] == 5'b10000 ? cell_80_7 :
    bitdata[600:596] == 5'b01000 ? cell_80_8 :
    bitdata[600:596] == 5'b11000 ? cell_80_9 :
    bitdata[600:596] == 5'b00100 ? cell_80_10 :
    bitdata[600:596] == 5'b10100 ? cell_80_11 :
    bitdata[600:596] == 5'b01100 ? cell_80_12 :
    bitdata[600:596] == 5'b11100 ? cell_80_13 :
    bitdata[600:596] == 5'b00010 ? cell_80_14 :
    bitdata[600:596] == 5'b10010 ? cell_80_15 :
    bitdata[600:596] == 5'b01010 ? cell_81_10 :
    bitdata[600:596] == 5'b11010 ? cell_81_11 :
    bitdata[600:596] == 5'b00110 ? cell_81_12 :
    bitdata[600:596] == 5'b10110 ? cell_81_13 :
    bitdata[600:596] == 5'b01110 ? cell_81_14 :
    bitdata[600:596] == 5'b11110 ? cell_81_15 :
    bitdata[600:596] == 5'b00001 ? cell_81_16 :
    bitdata[600:596] == 5'b10001 ? cell_81_17 :
    bitdata[600:596] == 5'b01001 ? cell_81_18 :
    bitdata[600:596] == 5'b11001 ? cell_81_19 :
    bitdata[600:596] == 5'b00101 ? cell_81_20 :
    bitdata[600:596] == 5'b10101 ? cell_81_21 :
    bitdata[600:596] == 5'b01101 ? cell_81_22 :
    bitdata[600:596] == 5'b11101 ? cell_81_23 :
    bitdata[600:596] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up5 =
   (bitdata[605:601] == 5'b00000 ? cell_80_6 :
    bitdata[605:601] == 5'b10000 ? cell_80_7 :
    bitdata[605:601] == 5'b01000 ? cell_80_8 :
    bitdata[605:601] == 5'b11000 ? cell_80_9 :
    bitdata[605:601] == 5'b00100 ? cell_80_10 :
    bitdata[605:601] == 5'b10100 ? cell_80_11 :
    bitdata[605:601] == 5'b01100 ? cell_80_12 :
    bitdata[605:601] == 5'b11100 ? cell_80_13 :
    bitdata[605:601] == 5'b00010 ? cell_80_14 :
    bitdata[605:601] == 5'b10010 ? cell_80_15 :
    bitdata[605:601] == 5'b01010 ? cell_81_10 :
    bitdata[605:601] == 5'b11010 ? cell_81_11 :
    bitdata[605:601] == 5'b00110 ? cell_81_12 :
    bitdata[605:601] == 5'b10110 ? cell_81_13 :
    bitdata[605:601] == 5'b01110 ? cell_81_14 :
    bitdata[605:601] == 5'b11110 ? cell_81_15 :
    bitdata[605:601] == 5'b00001 ? cell_81_16 :
    bitdata[605:601] == 5'b10001 ? cell_81_17 :
    bitdata[605:601] == 5'b01001 ? cell_81_18 :
    bitdata[605:601] == 5'b11001 ? cell_81_19 :
    bitdata[605:601] == 5'b00101 ? cell_81_20 :
    bitdata[605:601] == 5'b10101 ? cell_81_21 :
    bitdata[605:601] == 5'b01101 ? cell_81_22 :
    bitdata[605:601] == 5'b11101 ? cell_81_23 :
    bitdata[605:601] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up6 =
   (bitdata[610:606] == 5'b00000 ? cell_80_6 :
    bitdata[610:606] == 5'b10000 ? cell_80_7 :
    bitdata[610:606] == 5'b01000 ? cell_80_8 :
    bitdata[610:606] == 5'b11000 ? cell_80_9 :
    bitdata[610:606] == 5'b00100 ? cell_80_10 :
    bitdata[610:606] == 5'b10100 ? cell_80_11 :
    bitdata[610:606] == 5'b01100 ? cell_80_12 :
    bitdata[610:606] == 5'b11100 ? cell_80_13 :
    bitdata[610:606] == 5'b00010 ? cell_80_14 :
    bitdata[610:606] == 5'b10010 ? cell_80_15 :
    bitdata[610:606] == 5'b01010 ? cell_81_10 :
    bitdata[610:606] == 5'b11010 ? cell_81_11 :
    bitdata[610:606] == 5'b00110 ? cell_81_12 :
    bitdata[610:606] == 5'b10110 ? cell_81_13 :
    bitdata[610:606] == 5'b01110 ? cell_81_14 :
    bitdata[610:606] == 5'b11110 ? cell_81_15 :
    bitdata[610:606] == 5'b00001 ? cell_81_16 :
    bitdata[610:606] == 5'b10001 ? cell_81_17 :
    bitdata[610:606] == 5'b01001 ? cell_81_18 :
    bitdata[610:606] == 5'b11001 ? cell_81_19 :
    bitdata[610:606] == 5'b00101 ? cell_81_20 :
    bitdata[610:606] == 5'b10101 ? cell_81_21 :
    bitdata[610:606] == 5'b01101 ? cell_81_22 :
    bitdata[610:606] == 5'b11101 ? cell_81_23 :
    bitdata[610:606] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up7 =
   (bitdata[615:611] == 5'b00000 ? cell_80_6 :
    bitdata[615:611] == 5'b10000 ? cell_80_7 :
    bitdata[615:611] == 5'b01000 ? cell_80_8 :
    bitdata[615:611] == 5'b11000 ? cell_80_9 :
    bitdata[615:611] == 5'b00100 ? cell_80_10 :
    bitdata[615:611] == 5'b10100 ? cell_80_11 :
    bitdata[615:611] == 5'b01100 ? cell_80_12 :
    bitdata[615:611] == 5'b11100 ? cell_80_13 :
    bitdata[615:611] == 5'b00010 ? cell_80_14 :
    bitdata[615:611] == 5'b10010 ? cell_80_15 :
    bitdata[615:611] == 5'b01010 ? cell_81_10 :
    bitdata[615:611] == 5'b11010 ? cell_81_11 :
    bitdata[615:611] == 5'b00110 ? cell_81_12 :
    bitdata[615:611] == 5'b10110 ? cell_81_13 :
    bitdata[615:611] == 5'b01110 ? cell_81_14 :
    bitdata[615:611] == 5'b11110 ? cell_81_15 :
    bitdata[615:611] == 5'b00001 ? cell_81_16 :
    bitdata[615:611] == 5'b10001 ? cell_81_17 :
    bitdata[615:611] == 5'b01001 ? cell_81_18 :
    bitdata[615:611] == 5'b11001 ? cell_81_19 :
    bitdata[615:611] == 5'b00101 ? cell_81_20 :
    bitdata[615:611] == 5'b10101 ? cell_81_21 :
    bitdata[615:611] == 5'b01101 ? cell_81_22 :
    bitdata[615:611] == 5'b11101 ? cell_81_23 :
    bitdata[615:611] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up8 =
   (bitdata[620:616] == 5'b00000 ? cell_80_6 :
    bitdata[620:616] == 5'b10000 ? cell_80_7 :
    bitdata[620:616] == 5'b01000 ? cell_80_8 :
    bitdata[620:616] == 5'b11000 ? cell_80_9 :
    bitdata[620:616] == 5'b00100 ? cell_80_10 :
    bitdata[620:616] == 5'b10100 ? cell_80_11 :
    bitdata[620:616] == 5'b01100 ? cell_80_12 :
    bitdata[620:616] == 5'b11100 ? cell_80_13 :
    bitdata[620:616] == 5'b00010 ? cell_80_14 :
    bitdata[620:616] == 5'b10010 ? cell_80_15 :
    bitdata[620:616] == 5'b01010 ? cell_81_10 :
    bitdata[620:616] == 5'b11010 ? cell_81_11 :
    bitdata[620:616] == 5'b00110 ? cell_81_12 :
    bitdata[620:616] == 5'b10110 ? cell_81_13 :
    bitdata[620:616] == 5'b01110 ? cell_81_14 :
    bitdata[620:616] == 5'b11110 ? cell_81_15 :
    bitdata[620:616] == 5'b00001 ? cell_81_16 :
    bitdata[620:616] == 5'b10001 ? cell_81_17 :
    bitdata[620:616] == 5'b01001 ? cell_81_18 :
    bitdata[620:616] == 5'b11001 ? cell_81_19 :
    bitdata[620:616] == 5'b00101 ? cell_81_20 :
    bitdata[620:616] == 5'b10101 ? cell_81_21 :
    bitdata[620:616] == 5'b01101 ? cell_81_22 :
    bitdata[620:616] == 5'b11101 ? cell_81_23 :
    bitdata[620:616] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_8_up9 =
   (bitdata[625:621] == 5'b00000 ? cell_80_6 :
    bitdata[625:621] == 5'b10000 ? cell_80_7 :
    bitdata[625:621] == 5'b01000 ? cell_80_8 :
    bitdata[625:621] == 5'b11000 ? cell_80_9 :
    bitdata[625:621] == 5'b00100 ? cell_80_10 :
    bitdata[625:621] == 5'b10100 ? cell_80_11 :
    bitdata[625:621] == 5'b01100 ? cell_80_12 :
    bitdata[625:621] == 5'b11100 ? cell_80_13 :
    bitdata[625:621] == 5'b00010 ? cell_80_14 :
    bitdata[625:621] == 5'b10010 ? cell_80_15 :
    bitdata[625:621] == 5'b01010 ? cell_81_10 :
    bitdata[625:621] == 5'b11010 ? cell_81_11 :
    bitdata[625:621] == 5'b00110 ? cell_81_12 :
    bitdata[625:621] == 5'b10110 ? cell_81_13 :
    bitdata[625:621] == 5'b01110 ? cell_81_14 :
    bitdata[625:621] == 5'b11110 ? cell_81_15 :
    bitdata[625:621] == 5'b00001 ? cell_81_16 :
    bitdata[625:621] == 5'b10001 ? cell_81_17 :
    bitdata[625:621] == 5'b01001 ? cell_81_18 :
    bitdata[625:621] == 5'b11001 ? cell_81_19 :
    bitdata[625:621] == 5'b00101 ? cell_81_20 :
    bitdata[625:621] == 5'b10101 ? cell_81_21 :
    bitdata[625:621] == 5'b01101 ? cell_81_22 :
    bitdata[625:621] == 5'b11101 ? cell_81_23 :
    bitdata[625:621] == 5'b00011 ? cell_81_24 : 1'bx);
assign sw_0_1_9_down0 =
   (bitdata[464:460] == 5'b10001 ? sw_0_1_3_down0 :
    bitdata[464:460] == 5'b01001 ? sw_0_1_3_down1 :
    bitdata[464:460] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[464:460] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[464:460] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[464:460] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[464:460] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[464:460] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[464:460] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[464:460] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[464:460] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[464:460] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[464:460] == 5'b01010 ? sw_0_1_10_up0 :
    bitdata[464:460] == 5'b11010 ? sw_0_1_10_up1 :
    bitdata[464:460] == 5'b00110 ? sw_0_1_10_up2 :
    bitdata[464:460] == 5'b10110 ? sw_0_1_11_up0 :
    bitdata[464:460] == 5'b01110 ? sw_0_1_11_up1 :
    bitdata[464:460] == 5'b11110 ? sw_0_1_11_up2 :
    bitdata[464:460] == 5'b00001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_9_down1 =
   (bitdata[469:465] == 5'b10001 ? sw_0_1_3_down0 :
    bitdata[469:465] == 5'b01001 ? sw_0_1_3_down1 :
    bitdata[469:465] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[469:465] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[469:465] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[469:465] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[469:465] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[469:465] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[469:465] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[469:465] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[469:465] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[469:465] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[469:465] == 5'b01010 ? sw_0_1_10_up0 :
    bitdata[469:465] == 5'b11010 ? sw_0_1_10_up1 :
    bitdata[469:465] == 5'b00110 ? sw_0_1_10_up2 :
    bitdata[469:465] == 5'b10110 ? sw_0_1_11_up0 :
    bitdata[469:465] == 5'b01110 ? sw_0_1_11_up1 :
    bitdata[469:465] == 5'b11110 ? sw_0_1_11_up2 :
    bitdata[469:465] == 5'b00001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_9_down2 =
   (bitdata[474:470] == 5'b10001 ? sw_0_1_3_down0 :
    bitdata[474:470] == 5'b01001 ? sw_0_1_3_down1 :
    bitdata[474:470] == 5'b00000 ? sw_0_1_8_up0 :
    bitdata[474:470] == 5'b10000 ? sw_0_1_8_up1 :
    bitdata[474:470] == 5'b01000 ? sw_0_1_8_up2 :
    bitdata[474:470] == 5'b11000 ? sw_0_1_8_up3 :
    bitdata[474:470] == 5'b00100 ? sw_0_1_8_up4 :
    bitdata[474:470] == 5'b10100 ? sw_0_1_8_up5 :
    bitdata[474:470] == 5'b01100 ? sw_0_1_8_up6 :
    bitdata[474:470] == 5'b11100 ? sw_0_1_8_up7 :
    bitdata[474:470] == 5'b00010 ? sw_0_1_8_up8 :
    bitdata[474:470] == 5'b10010 ? sw_0_1_8_up9 :
    bitdata[474:470] == 5'b01010 ? sw_0_1_10_up0 :
    bitdata[474:470] == 5'b11010 ? sw_0_1_10_up1 :
    bitdata[474:470] == 5'b00110 ? sw_0_1_10_up2 :
    bitdata[474:470] == 5'b10110 ? sw_0_1_11_up0 :
    bitdata[474:470] == 5'b01110 ? sw_0_1_11_up1 :
    bitdata[474:470] == 5'b11110 ? sw_0_1_11_up2 :
    bitdata[474:470] == 5'b00001 ? sw_0_1_11_up3 : 1'bx);
assign sw_0_1_9_up0 = cell_43_0;
assign sw_1_0_1_down0 = sw_1_0_2_up0;
assign sw_1_0_1_up0 =
   (bitdata[912:911] == 2'b00 ? sw_1_0_3_up0 :
    bitdata[912:911] == 2'b10 ? sw_1_0_4_up0 :
    bitdata[912:911] == 2'b01 ? sw_1_0_4_up1 :
    bitdata[912:911] == 2'b11 ? sw_1_0_5_up0 : 8'bx);
assign sw_1_0_2_down0 = sw_1_0_1_up0;
assign sw_1_0_2_up0 =
   (bitdata[921:921] == 1'b0 ? sw_1_0_6_up0 :
    bitdata[921:921] == 1'b1 ? sw_1_0_7_up0 : 8'bx);
assign sw_1_0_3_down0 =
   (bitdata[914:913] == 2'b11 ? sw_1_0_1_down0 :
    bitdata[914:913] == 2'b00 ? sw_1_0_4_up0 :
    bitdata[914:913] == 2'b10 ? sw_1_0_4_up1 :
    bitdata[914:913] == 2'b01 ? sw_1_0_5_up0 : 8'bx);
assign sw_1_0_3_down1 =
   (bitdata[916:915] == 2'b11 ? sw_1_0_1_down0 :
    bitdata[916:915] == 2'b00 ? sw_1_0_4_up0 :
    bitdata[916:915] == 2'b10 ? sw_1_0_4_up1 :
    bitdata[916:915] == 2'b01 ? sw_1_0_5_up0 : 8'bx);
assign sw_1_0_3_up0 =
   (bitdata[924:923] == 2'b00 ? cell_73_7 :
    bitdata[924:923] == 2'b10 ? cell_87_0 :
    bitdata[924:923] == 2'b01 ? cell_89_0 : 8'bx);
assign sw_1_0_4_down0 =
   (bitdata[918:917] == 2'b01 ? sw_1_0_1_down0 :
    bitdata[918:917] == 2'b00 ? sw_1_0_3_up0 :
    bitdata[918:917] == 2'b10 ? sw_1_0_5_up0 : 8'bx);
assign sw_1_0_4_up0 =
   (bitdata[941:940] == 2'b00 ? cell_74_3 :
    bitdata[941:940] == 2'b10 ? cell_84_0 :
    bitdata[941:940] == 2'b01 ? cell_85_0 : 8'bx);
assign sw_1_0_4_up1 =
   (bitdata[943:942] == 2'b00 ? cell_74_3 :
    bitdata[943:942] == 2'b10 ? cell_84_0 :
    bitdata[943:942] == 2'b01 ? cell_85_0 : 8'bx);
assign sw_1_0_5_down0 =
   (bitdata[920:919] == 2'b11 ? sw_1_0_1_down0 :
    bitdata[920:919] == 2'b00 ? sw_1_0_3_up0 :
    bitdata[920:919] == 2'b10 ? sw_1_0_4_up0 :
    bitdata[920:919] == 2'b01 ? sw_1_0_4_up1 : 8'bx);
assign sw_1_0_5_up0 =
   (bitdata[951:951] == 1'b0 ? cell_75_3 :
    bitdata[951:951] == 1'b1 ? cell_86_0 : 8'bx);
assign sw_1_0_6_down0 =
   (bitdata[922:922] == 1'b1 ? sw_1_0_2_down0 :
    bitdata[922:922] == 1'b0 ? sw_1_0_7_up0 : 8'bx);
assign sw_1_0_6_up0 =
   (bitdata[958:958] == 1'b0 ? cell_69_1 :
    bitdata[958:958] == 1'b1 ? cell_70_1 : 8'bx);
assign sw_1_0_7_up0 =
   (bitdata[972:971] == 2'b00 ? cell_5_0 :
    bitdata[972:971] == 2'b10 ? cell_38_0 :
    bitdata[972:971] == 2'b01 ? cell_88_0 : 8'bx);
assign sw_1_1_1_down0 = sw_1_1_2_up0;
assign sw_1_1_1_up0 =
   (bitdata[974:973] == 2'b00 ? sw_1_1_3_up0 :
    bitdata[974:973] == 2'b10 ? sw_1_1_4_up0 :
    bitdata[974:973] == 2'b01 ? sw_1_1_4_up1 :
    bitdata[974:973] == 2'b11 ? sw_1_1_5_up0 : 8'bx);
assign sw_1_1_2_down0 = sw_1_1_1_up0;
assign sw_1_1_2_up0 = sw_1_1_6_up0;
assign sw_1_1_3_down0 =
   (bitdata[976:975] == 2'b11 ? sw_1_1_1_down0 :
    bitdata[976:975] == 2'b00 ? sw_1_1_4_up0 :
    bitdata[976:975] == 2'b10 ? sw_1_1_4_up1 :
    bitdata[976:975] == 2'b01 ? sw_1_1_5_up0 : 8'bx);
assign sw_1_1_3_up0 =
   (bitdata[985:984] == 2'b00 ? cell_74_3 :
    bitdata[985:984] == 2'b10 ? cell_86_0 :
    bitdata[985:984] == 2'b01 ? cell_87_0 :
    bitdata[985:984] == 2'b11 ? cell_89_0 : 8'bx);
assign sw_1_1_4_down0 =
   (bitdata[978:977] == 2'b01 ? sw_1_1_1_down0 :
    bitdata[978:977] == 2'b00 ? sw_1_1_3_up0 :
    bitdata[978:977] == 2'b10 ? sw_1_1_5_up0 : 8'bx);
assign sw_1_1_4_up0 =
   (bitdata[992:992] == 1'b0 ? cell_84_0 :
    bitdata[992:992] == 1'b1 ? cell_85_0 : 8'bx);
assign sw_1_1_4_up1 =
   (bitdata[993:993] == 1'b0 ? cell_84_0 :
    bitdata[993:993] == 1'b1 ? cell_85_0 : 8'bx);
assign sw_1_1_5_down0 =
   (bitdata[980:979] == 2'b11 ? sw_1_1_1_down0 :
    bitdata[980:979] == 2'b00 ? sw_1_1_3_up0 :
    bitdata[980:979] == 2'b10 ? sw_1_1_4_up0 :
    bitdata[980:979] == 2'b01 ? sw_1_1_4_up1 : 8'bx);
assign sw_1_1_5_down1 =
   (bitdata[982:981] == 2'b11 ? sw_1_1_1_down0 :
    bitdata[982:981] == 2'b00 ? sw_1_1_3_up0 :
    bitdata[982:981] == 2'b10 ? sw_1_1_4_up0 :
    bitdata[982:981] == 2'b01 ? sw_1_1_4_up1 : 8'bx);
assign sw_1_1_5_up0 =
   (bitdata[1003:1002] == 2'b00 ? cell_73_7 :
    bitdata[1003:1002] == 2'b10 ? cell_75_3 :
    bitdata[1003:1002] == 2'b01 ? cell_88_0 : 8'bx);
assign sw_1_1_6_down0 = sw_1_1_2_down0;
assign sw_1_1_6_up0 =
   (bitdata[1023:1022] == 2'b00 ? cell_5_0 :
    bitdata[1023:1022] == 2'b10 ? cell_38_0 :
    bitdata[1023:1022] == 2'b01 ? cell_69_1 :
    bitdata[1023:1022] == 2'b11 ? cell_70_1 : 8'bx);
assign sw_1_1_7_down0 =
   (bitdata[983:983] == 1'b1 ? sw_1_1_2_down0 :
    bitdata[983:983] == 1'b0 ? sw_1_1_6_up0 : 8'bx);
assign sw_2_0_1_down0 = sw_2_0_2_up0;
assign sw_2_0_1_up0 =
   (bitdata[1034:1033] == 2'b00 ? sw_2_0_3_up0 :
    bitdata[1034:1033] == 2'b10 ? sw_2_0_4_up0 :
    bitdata[1034:1033] == 2'b01 ? sw_2_0_5_up0 : 16'bx);
assign sw_2_0_2_down0 = sw_2_0_1_up0;
assign sw_2_0_2_up0 =
   (bitdata[1042:1041] == 2'b00 ? sw_2_0_6_up0 :
    bitdata[1042:1041] == 2'b10 ? sw_2_0_7_up0 :
    bitdata[1042:1041] == 2'b01 ? sw_2_0_8_up0 : 16'bx);
assign sw_2_0_3_down0 =
   (bitdata[1036:1035] == 2'b01 ? sw_2_0_1_down0 :
    bitdata[1036:1035] == 2'b00 ? sw_2_0_4_up0 :
    bitdata[1036:1035] == 2'b10 ? sw_2_0_5_up0 : 16'bx);
assign sw_2_0_3_up0 =
   (bitdata[1051:1049] == 3'b000 ? cell_62_5 :
    bitdata[1051:1049] == 3'b100 ? cell_63_6 :
    bitdata[1051:1049] == 3'b010 ? cell_63_7 :
    bitdata[1051:1049] == 3'b110 ? cell_93_0 :
    bitdata[1051:1049] == 3'b001 ? cell_94_0 : 16'bx);
assign sw_2_0_4_down0 =
   (bitdata[1038:1037] == 2'b01 ? sw_2_0_1_down0 :
    bitdata[1038:1037] == 2'b00 ? sw_2_0_3_up0 :
    bitdata[1038:1037] == 2'b10 ? sw_2_0_5_up0 : 16'bx);
assign sw_2_0_4_up0 =
   (bitdata[1062:1061] == 2'b00 ? cell_61_5 :
    bitdata[1062:1061] == 2'b10 ? cell_79_3 :
    bitdata[1062:1061] == 2'b01 ? cell_91_0 : 16'bx);
assign sw_2_0_5_down0 =
   (bitdata[1040:1039] == 2'b01 ? sw_2_0_1_down0 :
    bitdata[1040:1039] == 2'b00 ? sw_2_0_3_up0 :
    bitdata[1040:1039] == 2'b10 ? sw_2_0_4_up0 : 16'bx);
assign sw_2_0_5_up0 =
   (bitdata[1073:1072] == 2'b00 ? cell_67_1 :
    bitdata[1073:1072] == 2'b10 ? cell_72_3 :
    bitdata[1073:1072] == 2'b01 ? cell_77_2 :
    bitdata[1073:1072] == 2'b11 ? cell_78_3 : 16'bx);
assign sw_2_0_6_down0 =
   (bitdata[1044:1043] == 2'b01 ? sw_2_0_2_down0 :
    bitdata[1044:1043] == 2'b00 ? sw_2_0_7_up0 :
    bitdata[1044:1043] == 2'b10 ? sw_2_0_8_up0 : 16'bx);
assign sw_2_0_6_up0 =
   (bitdata[1091:1089] == 3'b000 ? cell_64_6 :
    bitdata[1091:1089] == 3'b100 ? cell_64_7 :
    bitdata[1091:1089] == 3'b010 ? cell_76_2 :
    bitdata[1091:1089] == 3'b110 ? cell_92_0 :
    bitdata[1091:1089] == 3'b001 ? cell_95_0 : 16'bx);
assign sw_2_0_7_down0 =
   (bitdata[1046:1045] == 2'b01 ? sw_2_0_2_down0 :
    bitdata[1046:1045] == 2'b00 ? sw_2_0_6_up0 :
    bitdata[1046:1045] == 2'b10 ? sw_2_0_8_up0 : 16'bx);
assign sw_2_0_7_up0 =
   (bitdata[1099:1098] == 2'b00 ? cell_65_2 :
    bitdata[1099:1098] == 2'b10 ? cell_66_1 :
    bitdata[1099:1098] == 2'b01 ? cell_71_3 : 16'bx);
assign sw_2_0_8_down0 =
   (bitdata[1048:1047] == 2'b01 ? sw_2_0_2_down0 :
    bitdata[1048:1047] == 2'b00 ? sw_2_0_6_up0 :
    bitdata[1048:1047] == 2'b10 ? sw_2_0_7_up0 : 16'bx);
assign sw_2_0_8_up0 =
   (bitdata[1114:1113] == 2'b00 ? cell_2_0 :
    bitdata[1114:1113] == 2'b10 ? cell_68_1 :
    bitdata[1114:1113] == 2'b01 ? cell_90_0 : 16'bx);
assign sw_2_1_1_down0 = sw_2_1_2_up0;
assign sw_2_1_1_up0 =
   (bitdata[1118:1117] == 2'b00 ? sw_2_1_3_up0 :
    bitdata[1118:1117] == 2'b10 ? sw_2_1_4_up0 :
    bitdata[1118:1117] == 2'b01 ? sw_2_1_5_up0 : 16'bx);
assign sw_2_1_2_down0 = sw_2_1_1_up0;
assign sw_2_1_2_up0 =
   (bitdata[1126:1125] == 2'b00 ? sw_2_1_6_up0 :
    bitdata[1126:1125] == 2'b10 ? sw_2_1_6_up1 :
    bitdata[1126:1125] == 2'b01 ? sw_2_1_7_up0 :
    bitdata[1126:1125] == 2'b11 ? sw_2_1_8_up0 : 16'bx);
assign sw_2_1_3_down0 =
   (bitdata[1120:1119] == 2'b01 ? sw_2_1_1_down0 :
    bitdata[1120:1119] == 2'b00 ? sw_2_1_4_up0 :
    bitdata[1120:1119] == 2'b10 ? sw_2_1_5_up0 : 16'bx);
assign sw_2_1_3_up0 =
   (bitdata[1135:1135] == 1'b0 ? cell_94_0 :
    bitdata[1135:1135] == 1'b1 ? cell_95_0 : 16'bx);
assign sw_2_1_4_down0 =
   (bitdata[1122:1121] == 2'b01 ? sw_2_1_1_down0 :
    bitdata[1122:1121] == 2'b00 ? sw_2_1_3_up0 :
    bitdata[1122:1121] == 2'b10 ? sw_2_1_5_up0 : 16'bx);
assign sw_2_1_4_up0 =
   (bitdata[1141:1140] == 2'b00 ? cell_71_3 :
    bitdata[1141:1140] == 2'b10 ? cell_78_3 :
    bitdata[1141:1140] == 2'b01 ? cell_92_0 :
    bitdata[1141:1140] == 2'b11 ? cell_93_0 : 16'bx);
assign sw_2_1_5_down0 =
   (bitdata[1124:1123] == 2'b01 ? sw_2_1_1_down0 :
    bitdata[1124:1123] == 2'b00 ? sw_2_1_3_up0 :
    bitdata[1124:1123] == 2'b10 ? sw_2_1_4_up0 : 16'bx);
assign sw_2_1_5_up0 =
   (bitdata[1156:1154] == 3'b000 ? cell_63_6 :
    bitdata[1156:1154] == 3'b100 ? cell_63_7 :
    bitdata[1156:1154] == 3'b010 ? cell_79_3 :
    bitdata[1156:1154] == 3'b110 ? cell_90_0 :
    bitdata[1156:1154] == 3'b001 ? cell_91_0 : 16'bx);
assign sw_2_1_6_down0 =
   (bitdata[1128:1127] == 2'b01 ? sw_2_1_2_down0 :
    bitdata[1128:1127] == 2'b00 ? sw_2_1_7_up0 :
    bitdata[1128:1127] == 2'b10 ? sw_2_1_8_up0 : 16'bx);
assign sw_2_1_6_up0 =
   (bitdata[1170:1169] == 2'b00 ? cell_67_1 :
    bitdata[1170:1169] == 2'b10 ? cell_68_1 :
    bitdata[1170:1169] == 2'b01 ? cell_72_3 :
    bitdata[1170:1169] == 2'b11 ? cell_77_2 : 16'bx);
assign sw_2_1_6_up1 =
   (bitdata[1172:1171] == 2'b00 ? cell_67_1 :
    bitdata[1172:1171] == 2'b10 ? cell_68_1 :
    bitdata[1172:1171] == 2'b01 ? cell_72_3 :
    bitdata[1172:1171] == 2'b11 ? cell_77_2 : 16'bx);
assign sw_2_1_7_down0 =
   (bitdata[1130:1129] == 2'b11 ? sw_2_1_2_down0 :
    bitdata[1130:1129] == 2'b00 ? sw_2_1_6_up0 :
    bitdata[1130:1129] == 2'b10 ? sw_2_1_6_up1 :
    bitdata[1130:1129] == 2'b01 ? sw_2_1_8_up0 : 16'bx);
assign sw_2_1_7_down1 =
   (bitdata[1132:1131] == 2'b11 ? sw_2_1_2_down0 :
    bitdata[1132:1131] == 2'b00 ? sw_2_1_6_up0 :
    bitdata[1132:1131] == 2'b10 ? sw_2_1_6_up1 :
    bitdata[1132:1131] == 2'b01 ? sw_2_1_8_up0 : 16'bx);
assign sw_2_1_7_up0 =
   (bitdata[1186:1185] == 2'b00 ? cell_2_0 :
    bitdata[1186:1185] == 2'b10 ? cell_65_2 :
    bitdata[1186:1185] == 2'b01 ? cell_66_1 :
    bitdata[1186:1185] == 2'b11 ? cell_76_2 : 16'bx);
assign sw_2_1_8_down0 =
   (bitdata[1134:1133] == 2'b11 ? sw_2_1_2_down0 :
    bitdata[1134:1133] == 2'b00 ? sw_2_1_6_up0 :
    bitdata[1134:1133] == 2'b10 ? sw_2_1_6_up1 :
    bitdata[1134:1133] == 2'b01 ? sw_2_1_7_up0 : 16'bx);
assign sw_2_1_8_up0 =
   (bitdata[1197:1196] == 2'b00 ? cell_61_5 :
    bitdata[1197:1196] == 2'b10 ? cell_62_5 :
    bitdata[1197:1196] == 2'b01 ? cell_64_6 :
    bitdata[1197:1196] == 2'b11 ? cell_64_7 : 16'bx);

endmodule
