----------------------------------------------------------------------------------
-- Company:     TU Vienna
-- Engineer:    Georg Blemenschitz
-- 
-- Create Date: 17:41:00 12/02/2009 
-- Design Name: FIFO
-- Module Name: tb_FIFOSync 
-- Description: VHDL Test Bench for module: FIFOSyncTop
--
-- Revision: 
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
 
entity tb_FIFOSync is
end tb_FIFOSync;

