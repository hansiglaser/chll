  constant TRFSM1Length : integer := 1778;
  constant TRFSM1Cfg    : std_logic_vector(TRFSM1Length-1 downto 0) := "00001100000000100000000100000010000101001100000000001000011000110001100000000000000011100010001100000000010000100000010100100000110000000101000001000100000100000000101100001100101000001000000110000000100100000100000011111100000000000000000000011111100000000000000000000000000000000010000100000000100001000000000000000000010001000011101100001000000000000100000000011000000100100000000000100000100000000010100100001100000000000100001000000000101000000000100010000000000010100000000011000010100100000010000000010100000000010100101100101100010000000100100000001001000011001100001000000000100100000001000100100100010001000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000011111100000000000000000000000000000000000001000000000110010000010001000000000000000010000000001100010010010001000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000111111000000000000000000000000000000000001111110000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000";
