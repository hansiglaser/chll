--------------------------------------------------------------------------------
-- Company:        vienna university of technology
-- Engineer:       mario faschang
-- Create Date:    11:12:56 19/01/2010
-- Module Name:    tb_I2CBusMaster
-- Project Name:   i2c master controller
-- Description:  * testbench for I2CBusMaster
--               * generates different scenarios of the i2c-bus-communication
--                 to verify the behavior of the i2cBusMaster.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY tb_I2CBusMaster IS

END tb_I2CBusMaster;

