----------------------------------------------------------------------------------
-- Company:  TU Vienna
-- Engineer: Armin FALTINGER
--
-- Create Date:    13:46:24 11/21/2009
-- Project Name:   Uart
-- Module Name:    ErrorIndicator - structure
-- Dependencies:   Module to bind 3 instances of ErrorBit.vhd
--                   instances are PARITYERR, STOPERR and RXBUFFERR
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- if an error (Parity, Stopbit or RxBufferFull) occurs
--   the status is indicated on the output
-- the errors are cleared by a master reset or a ErrorReset just for the module
-- RxBufferFull error means that the Fifo is full, but data is still received

entity ErrorIndicator is
  Port ( -- Errors generated by the TX/RX module
         ParityError_i                : in   STD_LOGIC;
         StopBitError_i               : in   STD_LOGIC;
         RxBufferFullError_i          : in   STD_LOGIC;
         -- general inputs
         Clk_i                        : in   STD_LOGIC;
         Reset_i_n                    : in   STD_LOGIC;
         ErrorReset_i                 : in   STD_LOGIC;
         -- Indication
         StopBitErrorIndicator_o      : out  STD_LOGIC;
         ParityErrorIndicator_o       : out  STD_LOGIC;
         RxBufferFullErrorIndicator_o : out  STD_LOGIC
        );
end ErrorIndicator;

