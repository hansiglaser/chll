  constant bitdataLength : integer := 1282;
  constant bitdataCfg    : std_logic_vector(bitdataLength-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000010000000000000000000000000000000000000000001000000000000000000000000000000000010001000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000110010010010110001000001111010010000100000000000101011010010011110000001001111000000000000000000000000000000000000000000000000000000000000001000000110010100000000000000000000";
