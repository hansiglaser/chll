  constant SPIFSMLength : integer := 1295;
  constant SPIFSMCfg    : std_logic_vector(SPIFSMLength-1 downto 0) := "00001001010000000000010010001000110000000000000000000110000000000000001001000100000100000000001000000010100011000000000010010000000000000101000000000000000100000000000000001100010000000000010000000110000000100100001000000000001100001100000001010001100000000000000001111100000000000000000000000000000011111000000000000000000000000000000111110000000000000000000000000000001111100000000000000000000000000000011111000000000000000000000000000000111110000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
