  constant SPIFSMLength : integer := 1295;
  constant SPIFSMCfg    : std_logic_vector(SPIFSMLength-1 downto 0) := "00001001000000000000010100001000101000000000000000000110001000000000001000011111000000000000000000001111100000000000000000000000000000000101000000000000001000000000000000001100001100000000001000000100000000010100000000000000100001001000000000110000110000000000100010010100000010010000100000000000110000101000000101000101000000000000000111110000000000000000000000000000001111100000000000000000000000000000011111000000000000000000000000000000111110000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
