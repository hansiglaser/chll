  constant SPIFSMLength : integer := 1295;
  constant SPIFSMCfg    : std_logic_vector(SPIFSMLength-1 downto 0) := "00001001000000000001000000001000101000000000000010000110001000000000000010011111000000000000000000001111100000000000000000000000000000000101000000000000000010000000000000001100001100000000000100000100000000010100000000000000010000001000000000110000110000000000100000010100000010010000100000000000000100101000000101000101000000000000001111110000000000000000000000000000001111100000000000000000000000000000011111000000000000000000000000000000111110000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
