  constant ReconfSignalsLength : integer := 9;
  constant ReconfSignalsCfg    : std_logic_vector(ReconfSignalsLength-1 downto 0) := "000000000";
