-- Automatically generated: write_netlist -wrapapp -vhdl -instance reconflogic-wrapslowadt7410-instance.vhd

  MyReconfigLogic_0: MyReconfigLogic
    port map (
      Reset_n_i => Reset_n_s,
      Clk_i => Clk_i,
      AdcConvComplete_i => AdcConvComplete_i,
      AdcDoConvert_o => AdcDoConvert_o,
      AdcValue_i => AdcValue_i,
      I2C_Busy_i => I2C_Busy,
      I2C_DataIn_o => I2C_DataIn,
      I2C_DataOut_i => I2C_DataOut,
      I2C_Divider800_o => I2C_Divider800,
      I2C_ErrAckParam_o => I2C_ErrAckParam,
      I2C_Error_i => I2C_Error,
      I2C_F100_400_n_o => I2C_F100_400_n,
      I2C_FIFOEmpty_i => I2C_FIFOEmpty,
      I2C_FIFOFull_i => I2C_FIFOFull,
      I2C_FIFOReadNext_o => I2C_FIFOReadNext,
      I2C_FIFOWrite_o => I2C_FIFOWrite,
      I2C_ReadCount_o => I2C_ReadCount,
      I2C_ReceiveSend_n_o => I2C_ReceiveSend_n,
      I2C_StartProcess_o => I2C_StartProcess,
      Inputs_i => Inputs_i,
      Outputs_o => Outputs_o,
      ReconfModuleIRQs_o => ReconfModuleIRQs_s,
      SPI_CPHA_o => SPI_CPHA,
      SPI_CPOL_o => SPI_CPOL,
      SPI_DataIn_o => SPI_DataIn,
      SPI_DataOut_i => SPI_DataOut,
      SPI_FIFOEmpty_i => SPI_FIFOEmpty,
      SPI_FIFOFull_i => SPI_FIFOFull,
      SPI_LSBFE_o => SPI_LSBFE,
      SPI_ReadNext_o => SPI_ReadNext,
      SPI_SPPR_SPR_o => SPI_SPPR_SPR,
      SPI_Transmission_i => SPI_Transmission,
      SPI_Write_o => SPI_Write,
      ReconfModuleIn_i => ReconfModuleIn_s,
      ReconfModuleOut_o => ReconfModuleOut_s,
      I2C_Errors_i => I2C_Errors,
      PerAddr_i => Per_Addr_s,
      PerDIn_i => Per_DIn_s,
      PerWr_i => Per_Wr_s,
      PerEn_i => Per_En_s,
      CfgIntfDOut_o => CfgIntf_DOut_s,
      ParamIntfDOut_o => ParamIntf_DOut_s
    );

