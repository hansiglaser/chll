  constant SPIFSMLength : integer := 1295;
  constant SPIFSMCfg    : std_logic_vector(SPIFSMLength-1 downto 0) := "00001001110000100110010000010000000000000111000000001010101000000100101000000110000110000010010000100011100100000010011000100000000000010001000000000001110000000000000000100100011000000100100000000010000000010100010000000010100001000100000000110010000000010010000010001100000010100001100000000100000000011000000100101001000010001000000010000000000011001010000010010100000100100000000110001000001000010000001010000000100100001000010001000000010100000001010010100000000010000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000111110000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000";
